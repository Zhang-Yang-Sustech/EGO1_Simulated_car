`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/01/05 19:55:32
// Design Name: 
// Module Name: Vga
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module vga_control(
input wire vga_clk,
input wire sys_rst,
input wire [11:0] pix_data,//��ĳ���������Ϣ
output reg [9:0] pix_x,
output reg [9:0] pix_y,
output wire[0:0] hsync,
output wire[0:0] vsync,
output reg [11:0] vga_rgb
);

parameter H_SYNC =10'd96; //��ͬ������
parameter H_BA=10'd48;
parameter H_VA = 10'd640; //�Ϸ���ʾ����
parameter H_TO=10'd800;

parameter V_SYNC =10'd2; //��ͬ������
parameter V_BA=10'd33;
parameter V_VA = 10'd480; //�Ϸ���ʾ����
parameter V_TO=10'd525;

reg[9:0] cnt_h=10'b00000_00001;
reg[9:0] cnt_v=10'b00000_00001;


    
        always@(posedge vga_clk,posedge sys_rst)begin
        if(sys_rst==1'b1)begin
            cnt_v<=10'b00000_00001;
            end
            else if( (cnt_h==H_TO)&& (cnt_v < V_TO  ) ) begin
                cnt_v<=cnt_v+10'b00000_00001;
            end
            else if( (cnt_h ==H_TO) &&(cnt_v == V_TO  )  ) begin
                cnt_v<=10'b00000_00001;
            end
            else begin
            cnt_v <=cnt_v;
            end
        end
        
        always@(posedge vga_clk,posedge sys_rst)begin
             if(sys_rst==1'b1)begin
       cnt_h<=0;
       end
       else if(cnt_h ==(H_TO) ) begin
           cnt_h<=10'b00000_00001;
       end
       else begin
       cnt_h<=cnt_h+10'b00000_00001;
       end
        end



           always@(posedge  vga_clk)begin
                  if( (cnt_h >=H_SYNC +H_BA-1'b1)&& (cnt_h <H_SYNC +H_BA + H_VA-1'b1) &&
                     (cnt_v >= V_SYNC +V_BA ) && (cnt_v <V_SYNC +V_BA + V_VA)  )begin
                        pix_x <=cnt_h -(H_SYNC +H_BA ) ;
                        pix_y <=cnt_v-(V_SYNC +V_BA );
                    end
                    else begin
                        pix_x<=10'b00000_00000;
                        pix_y<=10'b00000_00000;
                    end
            end
            
                always@(posedge  vga_clk)begin
                          if( (cnt_h >=H_SYNC +H_BA)&& (cnt_h <H_SYNC +H_BA + H_VA) &&
                             (cnt_v >= V_SYNC +V_BA ) && (cnt_v <V_SYNC +V_BA + V_VA)  )begin
                              vga_rgb<=pix_data;
                            end
                            else begin
                                vga_rgb<=12'b0000_0000_0000;
                            end
                    end
            
            assign hsync =(cnt_h <=H_SYNC  ? 1'b0:1'b1);
            assign vsync =(cnt_v <= V_SYNC  ? 1'b0 :1'b1);
            
 endmodule

module vga_draw(//25MHz
input wire vga_clk,
input wire sys_rst,
input wire [3:0]state,
input wire [2:0]swi,

input wire [9:0]pix_x,
input wire [9:0]pix_y,
output reg [11:0] pix_data
);
parameter off =4'b0000, no_st = 4'b0011, start = 4'b0111, movef = 4'b0110, moveb = 4'b0101;
//�ֶ�ģʽ���״̬���ֱ�Ϊ�ػ���δ�𲽡��𲽡�ǰ�������ˣ��ɿ������ҷ���
parameter wait_command=4'b1000,left_turning=4'b1001,right_turning=4'b1010,circle_turning=4'b1011,keep_go=4'b1110,semi_movef=4'b1111;
//�ֱ�Ϊ�ȴ�ָ���ת����ת����ͷ������ǰ�������ɿ������ҷ����ǰ��
parameter black = 12'h000, blue = 12'h00f, white = 12'hfff;
reg [255:0] char0 [63:0];
reg [255:0] char1 [63:0];
reg [255:0] char2 [63:0];
reg [255:0] char00 [63:0];//�ֶ�
reg [255:0] char00_1 [63:0];//���Զ�
reg [255:0] char00_2 [63:0];//ȫ�Զ�
reg [255:0] char11 [63:0];//�ػ�
reg [255:0] char11_1 [63:0];//δ��
reg [255:0] char11_2 [63:0];//��
reg [255:0] char11_3 [63:0];//�ƶ�
reg [255:0] char11_4 [63:0];//�ȴ�ָ��
reg [255:0] char11_5 [63:0];//ת��
reg [255:0] char11_6 [63:0];//��ͷ
reg [31:0] char22_0 [63:0];//0
reg [31:0] char22_1 [63:0];//1
reg [31:0] char22_2 [63:0];//2
reg [31:0] char22_3 [63:0];//3
reg [127:0] char22_4 [63:0];//4
//reg [95:0] char22_5 [63:0];//5

reg [511:0] char   [479:0];
parameter onekm = 37'd2500_0000,tenkm = 37'd25000_0000,hkm = 37'd250000_0000,diankm = 37'd250_0000;
reg[36:0] li;
always@(posedge vga_clk) begin
    case(state)
        off: li<=0;
        movef: li <= li+1'b1;
        moveb: li <= li+1'b1;
        semi_movef: li <= li+1'b1;
        keep_go: li <= li+1'b1;
        default: li <= li;
    endcase
end

always@(posedge vga_clk) begin
char0[  0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char0[  1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char0[  2] <= 256'h000E0000E00E0000000000000000000000000000000000000000000000000000;
char0[  3] <= 256'h000F8000F80F8000000000001000000000000000000000000000000000000000;
char0[  4] <= 256'h000FE000FE0FE000000000001C00000000000000000000000000000000000000;
char0[  5] <= 256'h000FE000FC0FC000000000001F00000000000000000000000000000000000000;
char0[  6] <= 256'h000F8000F80F8000000000001F0E000000000000000000000000000000000000;
char0[  7] <= 256'h000F8000F80F8180000000001E07800000000000000000000000000000000000;
char0[  8] <= 256'h000F8000F80F83C0000000001E03E00000000000000000000000000000000000;
char0[  9] <= 256'h000F8000F80F87E0000000001E01F00000000000000000000000000000000000;
char0[10] <= 256'h000F83FFFFFFFFF0000000001E00F80000000000000000000000000000000000;
char0[11] <= 256'h000F81FFFFFFFFF8000000001E00F80000000000000000000000000000000000;
char0[12] <= 256'h000F80C0F80F8000000000001E00780000000000000000000000000000000000;
char0[13] <= 256'h000F8000F80F8000000000001E007A0000000000000000000000000000000000;
char0[14] <= 256'h000F8600F80F8000000000001E00370000000000000000000000000000000000;
char0[15] <= 256'h000F8F00F80F8000000000001E000F8000000000000000000000000000000000;
char0[16] <= 256'h000F9F80F80F8000000000001E001FC000000000000000000000000000000000;
char0[17] <= 256'h3FFFFFC0F00E000007FFFFFFFFFFFFE000000000000000000000000000000000;
char0[18] <= 256'h1FFFFFE8C000180003FFFFFFFFFFFFF000000000000000000000000000000000;
char0[19] <= 256'h0C0F800E00003C00018000000E00000000000000000000000000000000000000;
char0[20] <= 256'h001F800FFFFFFE00000000000E00000000000000000000000000000000000000;
char0[21] <= 256'h001F800FFFFFFF00000000000E00000000000000000000000000000000000000;
char0[22] <= 256'h001F800F80007E00000000000E00000000000000000000000000000000000000;
char0[23] <= 256'h001F800F80007C00000000000E00000000000000000000000000000000000000;
char0[24] <= 256'h001F800F80007C00000000000F00000000000000000000000000000000000000;
char0[25] <= 256'h003FC00F80007C00000000000F00000000000000000000000000000000000000;
char0[26] <= 256'h003FF00F80007C00000000040F00000000000000000000000000000000000000;
char0[27] <= 256'h003FFC0FFFFFFC000000000E0F00000000000000000000000000000000000000;
char0[28] <= 256'h007FFE0FFFFFFC000000001F0F00000000000000000000000000000000000000;
char0[29] <= 256'h007FBF0F80007C0003FFFFFF8700000000000000000000000000000000000000;
char0[30] <= 256'h007F9F8F80007C0001FFFFFFC700000000000000000000000000000000000000;
char0[31] <= 256'h00FF9F8F80007C0000803C000780000000000000000000000000000000000000;
char0[32] <= 256'h00FF8F8F80007C0000003C0007800000001E0000000000000000000000000000;
char0[33] <= 256'h00FF8F8F80007C0000003C0007800000007F8000000000000000000000000000;
char0[34] <= 256'h01FF878F80007C0000003C0007800000007F8000000000000000000000000000;
char0[35] <= 256'h01EF878FFFFFFC0000003C000380000000FF8000000000000000000000000000;
char0[36] <= 256'h03CF830FFFFFFC0000003C0003C0000000FFC000000000000000000000000000;
char0[37] <= 256'h03CF800F87C07C0000003C0003C0000000FF8000000000000000000000000000;
char0[38] <= 256'h078F800F87C07C0000003C0003C00000007F8000000000000000000000000000;
char0[39] <= 256'h078F800F07C0780000003C0001E00000007F0000000000000000000000000000;
char0[40] <= 256'h0F0F800807C0000000003C0001E00000001C0000000000000000000000000000;
char0[41] <= 256'h0E0F800007C001C000003C0001F0000000000000000000000000000000000000;
char0[42] <= 256'h1E0F800007C003E000003C0000F0000000000000000000000000000000000000;
char0[43] <= 256'h1C0F800007C007F000003C0000F0002000000000000000000000000000000000;
char0[44] <= 256'h380F8FFFFFFFFFF800003C000078002000000000000000000000000000000000;
char0[45] <= 256'h300F8FFFFFFFFFFC00003C000078006000000000000000000000000000000000;
char0[46] <= 256'h000F87C00FF0000000003C00383C006000000000000000000000000000000000;
char0[47] <= 256'h000F80000FB8000000003C03E03E0060003E0000000000000000000000000000;
char0[48] <= 256'h000F80001F38000000003C7F001E0060007F0000000000000000000000000000;
char0[49] <= 256'h000F80001F1C000000003FF8001F006000FF8000000000000000000000000000;
char0[50] <= 256'h000F80003E1E000000007FC0000F806000FF8000000000000000000000000000;
char0[51] <= 256'h000F80007E0F00000007FE000007C0E000FF8000000000000000000000000000;
char0[52] <= 256'h000F80007C07C00000FFF0000007F0E000FF8000000000000000000000000000;
char0[53] <= 256'h000F8000F807E0000FFF80000003F8E0007F8000000000000000000000000000;
char0[54] <= 256'h000F8001F003F80007FC00000001FEE0007F0000000000000000000000000000;
char0[55] <= 256'h000F8003E001FF0007E000000000FFE0001C0000000000000000000000000000;
char0[56] <= 256'h000F8007C000FFF80380000000003FF000000000000000000000000000000000;
char0[57] <= 256'h000F801F80007FFC0100000000001FF000000000000000000000000000000000;
char0[58] <= 256'h000F807F00003FF000000000000007F000000000000000000000000000000000;
char0[59] <= 256'h000F81FC00000FC000000000000001F800000000000000000000000000000000;
char0[60] <= 256'h000F8FE000000380000000000000003800000000000000000000000000000000;
char0[61] <= 256'h000E3F0000000000000000000000000000000000000000000000000000000000;
char0[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char0[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;

   char1[  0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char1[  1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char1[  2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char1[  3] <= 256'h000070000C0000000000000C0000000000000000000000000000000000000000;
 char1[  4] <= 256'h00007C000F0000000000000F0000000000000000000000000000000000000000;
 char1[  5] <= 256'h00007F000FC000000000000FC000000000000000000000000000000000000000;
 char1[  6] <= 256'h00007E000FE600000000000FC000000000000000000000000000000000000000;
 char1[  7] <= 256'h00007C000FC780000000000F0000000000000000000000000000000000000000;
 char1[  8] <= 256'h00007C000F83E0000000000F0000000000000000000000000000000000000000;
 char1[  9] <= 256'h00007C000F81F8000000000F0000000000000000000000000000000000000000;
 char1[10] <= 256'h00007C000F80FE000000000F0000000000000000000000000000000000000000;
 char1[11] <= 256'h00007C000F80FE000000000F0000060000000000000000000000000000000000;
 char1[12] <= 256'h00007C000F807F000000000F00000F0000000000000000000000000000000000;
 char1[13] <= 256'h0C007C000F803F000000000E00001F8000000000000000000000000000000000;
 char1[14] <= 256'h0E007C000F803F000FFFFFFFFFFFFFC000000000000000000000000000000000;
 char1[15] <= 256'h0F007C000F801F0007FFFFFFFFFFFFE000000000000000000000000000000000;
 char1[16] <= 256'h07C07C000F801F000200001EC000000000000000000000000000000000000000;
 char1[17] <= 256'h03E07C000F800E000000001C4000000000000000000000000000000000000000;
 char1[18] <= 256'h03F07C000F8006000000003C6000000000000000000000000000000000000000;
 char1[19] <= 256'h01F87C000F8000000000003C3000000000000000000000000000000000000000;
 char1[20] <= 256'h01F87C000F800380000000383000000000000000000000000000000000000000;
 char1[21] <= 256'h00FC7C000F8007C0000000781800000000000000000000000000000000000000;
 char1[22] <= 256'h00FC7C000F800FE0000000700C00000000000000000000000000000000000000;
 char1[23] <= 256'h00FC7FFFFFFFFFF0000000F00E00000000000000000000000000000000000000;
 char1[24] <= 256'h007C7FFFFFFFFFF8000001E00700000000000000000000000000000000000000;
 char1[25] <= 256'h007C7DF00FF00000000001E00380000000000000000000000000000000000000;
 char1[26] <= 256'h00787C000FF00000000003C001C0000000000000000000000000000000000000;
 char1[27] <= 256'h00387C000FF000000000078001F0000000000000000000000000000000000000;
 char1[28] <= 256'h00007C001FF0000000000FC000F8000000000000000000000000000000000000;
 char1[29] <= 256'h00007C001F70000000001F78007E000000000000000000000000000000000000;
 char1[30] <= 256'h00007C001F78000000003C3E003F800000000000000000000000000000000000;
 char1[31] <= 256'h00007C001F3800000000781F001FE00000000000000000000000000000000000;
 char1[32] <= 256'h0000FC001F3800000001F00FC007FC00001E0000000000000000000000000000;
 char1[33] <= 256'h0001FC001F3800000003C007E003FFE0007F8000000000000000000000000000;
 char1[34] <= 256'h0003FC001F3C0000000F0003E000FFF8007F8000000000000000000000000000;
 char1[35] <= 256'h000FFC003F3C0000003C0001E0003FC000FF8000000000000000000000000000;
 char1[36] <= 256'h001F7C003E3C000000F00000E0000F0000FFC000000000000000000000000000;
 char1[37] <= 256'h003E7C003E1E000007800000E000030000FF8000000000000000000000000000;
 char1[38] <= 256'h007C7C003E1E00001C00003000000000007F8000000000000000000000000000;
 char1[39] <= 256'h01F87C003E1F00000000181C00000000007F0000000000000000000000000000;
 char1[40] <= 256'h03F07C007C0F000000001E0F00000000001C0000000000000000000000000000;
 char1[41] <= 256'h0FE07C007C0F000000001F878000000000000000000000000000000000000000;
 char1[42] <= 256'h3FC07C007C0F800000081E07E001800000000000000000000000000000000000;
 char1[43] <= 256'h3F807C00F80F800000081E03E000E00000000000000000000000000000000000;
 char1[44] <= 256'h1F807C00F807C00000181E01F000700000000000000000000000000000000000;
 char1[45] <= 256'h0F007C01F007C00000181E01F0007C0000000000000000000000000000000000;
 char1[46] <= 256'h0E007C01F003E00000381E00F0103E0000000000000000000000000000000000;
 char1[47] <= 256'h06007C01F003F00000381E00E0101F00003E0000000000000000000000000000;
 char1[48] <= 256'h00007C03E001F00000781E0040101F80007F0000000000000000000000000000;
 char1[49] <= 256'h00007C03C001F80000F81E0000100F8000FF8000000000000000000000000000;
 char1[50] <= 256'h00007C07C000FC0000F01E0000100F8000FF8000000000000000000000000000;
 char1[51] <= 256'h00007C0F8000FE0003F01E000018078000FF8000000000000000000000000000;
 char1[52] <= 256'h00007C0F80007F0007F01E000038078000FF8000000000000000000000000000;
 char1[53] <= 256'h00007C1F00007F8007E01C0000380300007F8000000000000000000000000000;
 char1[54] <= 256'h00007C3E00003FE007C01E00003C0000007F0000000000000000000000000000;
 char1[55] <= 256'h00007C3C00001FF000001E00007E0000001C0000000000000000000000000000;
 char1[56] <= 256'h00007C7800001FFC00001FFFFFFE000000000000000000000000000000000000;
 char1[57] <= 256'h00007CF000000FFC00000FFFFFFC000000000000000000000000000000000000;
 char1[58] <= 256'h00007DE0000007C0000007FFFFF8000000000000000000000000000000000000;
 char1[59] <= 256'h00007FC000000380000000000000000000000000000000000000000000000000;
 char1[60] <= 256'h0000778000000000000000000000000000000000000000000000000000000000;
 char1[61] <= 256'h00004E0000000000000000000000000000000000000000000000000000000000;
 char1[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char1[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    
 char2[  0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char2[  1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char2[  2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char2[  3] <= 256'h0000000000000000000001000000000000000000000000000000000000000000;
 char2[  4] <= 256'h0000000000000000000007820000020000000000000000000000000000000000;
 char2[  5] <= 256'h000600000001C00000001FC18000070000000000000000000000000000000000;
 char2[  6] <= 256'h000700000003E0000000FFC1FFFFFF8000000000000000000000000000000000;
 char2[  7] <= 256'h0007FFFFFFFFF0000007FFE1FFFFFFC000000000000000000000000000000000;
 char2[  8] <= 256'h0007FFFFFFFFF800007FF001C000078000000000000000000000000000000000;
 char2[  9] <= 256'h0007C007C003F00007FDC001C000070000000000000000000000000000000000;
 char2[10] <= 256'h0007C007C003E0000801C001C000070000000000000000000000000000000000;
 char2[11] <= 256'h0007C007C003E0000001C001C000070000000000000000000000000000000000;
 char2[12] <= 256'h0007C007C003E0000001C001C000070000000000000000000000000000000000;
 char2[13] <= 256'h0007C007C003E0000001C001C000070000000000000000000000000000000000;
 char2[14] <= 256'h0007C007C003E0000001C001C000070000000000000000000000000000000000;
 char2[15] <= 256'h0007C007C003E0000001C001C000070000000000000000000000000000000000;
 char2[16] <= 256'h0007C007C003E0000001C001C000070000000000000000000000000000000000;
 char2[17] <= 256'h0007C007C003E0000001C001C000070000000000000000000000000000000000;
 char2[18] <= 256'h0007C007C003E0000001C001C000070000000000000000000000000000000000;
 char2[19] <= 256'h0007FFFFFFFFE0000001C081C000070000000000000000000000000000000000;
 char2[20] <= 256'h0007FFFFFFFFE0000001C1C1C000070000000000000000000000000000000000;
 char2[21] <= 256'h0007C007C003E0003FFFFFE1FFFFFF0000000000000000000000000000000000;
 char2[22] <= 256'h0007C007C003E0001FFFFFF1FFFFFF0000000000000000000000000000000000;
 char2[23] <= 256'h0007C007C003E0000C03C001C000070000000000000000000000000000000000;
 char2[24] <= 256'h0007C007C003E0000003C001C000070000000000000000000000000000000000;
 char2[25] <= 256'h0007C007C003E0000007C001C000040000000000000000000000000000000000;
 char2[26] <= 256'h0007C007C003E0000007C0010000000000000000000000000000000000000000;
 char2[27] <= 256'h0007C007C003E0000007C0000000000000000000000000000000000000000000;
 char2[28] <= 256'h0007C007C003E0000007F0000000018000000000000000000000000000000000;
 char2[29] <= 256'h0007C007C003E000000FDC00000003C000000000000000000000000000000000;
 char2[30] <= 256'h0007C007C003E000000FCE1FFFFFFFE000000000000000000000000000000000;
 char2[31] <= 256'h0007C007C003E000000FC78FFFFFFFF000000000000000000000000000000000;
 char2[32] <= 256'h0007FFFFFFFFE000001FC7C600780000001E0000000000000000000000000000;
 char2[33] <= 256'h0007FFFFFFFFE000001DC3C000780000007F8000000000000000000000000000;
 char2[34] <= 256'h0007C007C003E000001DC3C000780000007F8000000000000000000000000000;
 char2[35] <= 256'h0007C007C003E0000039C1C00078000000FF8000000000000000000000000000;
 char2[36] <= 256'h0007C007C003C0000039C1C00078000000FFC000000000000000000000000000;
 char2[37] <= 256'h00070007C00000000071C0C00078000000FF8000000000000000000000000000;
 char2[38] <= 256'h00000007C00000000071C00000780000007F8000000000000000000000000000;
 char2[39] <= 256'h00000007C00000000061C00000780000007F0000000000000000000000000000;
 char2[40] <= 256'h00000007C000000000E1C00000780200001C0000000000000000000000000000;
 char2[41] <= 256'h00000007C000700000C1C0000078070000000000000000000000000000000000;
 char2[42] <= 256'h00000007C000F80001C1C007FFFFFF8000000000000000000000000000000000;
 char2[43] <= 256'h00000007C001FC000181C003FFFFFFC000000000000000000000000000000000;
 char2[44] <= 256'h00FFFFFFFFFFFE000301C0010078000000000000000000000000000000000000;
 char2[45] <= 256'h007FFFFFFFFFFF000301C0000078000000000000000000000000000000000000;
 char2[46] <= 256'h003E0007C00000000601C0000078000000000000000000000000000000000000;
 char2[47] <= 256'h00000007C00000000C01C00000780000003E0000000000000000000000000000;
 char2[48] <= 256'h00000007C00000000801C00000780000007F0000000000000000000000000000;
 char2[49] <= 256'h00000007C00000001801C0000078000000FF8000000000000000000000000000;
 char2[50] <= 256'h00000007C00000003001C0000078000000FF8000000000000000000000000000;
 char2[51] <= 256'h00000007C00000000001C0000078000000FF8000000000000000000000000000;
 char2[52] <= 256'h00000007C00000000001C0000078004000FF8000000000000000000000000000;
 char2[53] <= 256'h00000007C00001800001C000007800C0007F8000000000000000000000000000;
 char2[54] <= 256'h00000007C00003C00001C000007801E0007F0000000000000000000000000000;
 char2[55] <= 256'h00000007C00007E00001C1FFFFFFFFF0001C0000000000000000000000000000;
 char2[56] <= 256'h00000007C0000FF00001C0FFFFFFFFF800000000000000000000000000000000;
 char2[57] <= 256'h1FFFFFFFFFFFFFF00001C0600000000000000000000000000000000000000000;
 char2[58] <= 256'h1FFFFFFFFFFFFFF80001C0000000000000000000000000000000000000000000;
 char2[59] <= 256'h0F800000000000000001C0000000000000000000000000000000000000000000;
 char2[60] <= 256'h0000000000000000000100000000000000000000000000000000000000000000;
 char2[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char2[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 char2[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 
 
 case(swi)
    3'b000: begin//�ػ�
             char00[  0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
             char00[  1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
             char00[  2] <= 256'h0000000000000000000200000000000000000000000000000000000000000000;
             char00[  3] <= 256'h0000600000E00000000380000000000000000000000000000000000000000000;
             char00[  4] <= 256'h0000780000F800000003E0000000000000000000000000000000000000000000;
             char00[  5] <= 256'h00003E0000FC00000003C0000000000000000000000000000000000000000000;
             char00[  6] <= 256'h00001F0001FF0000000380000000000000000000000000000000000000000000;
             char00[  7] <= 256'h00000F8001FE0000000380020001000000000000000000000000000000000000;
             char00[  8] <= 256'h00000FC001F80000000380038003800000000000000000000000000000000000;
             char00[  9] <= 256'h000007E003F0000000038003FFFFE00000000000000000000000000000000000;
             char00[10] <= 256'h000003F003E0000000038003FFFFF00000000000000000000000000000000000;
             char00[11] <= 256'h000003F803E0000000038003C003C00000000000000000000000000000000000;
             char00[12] <= 256'h000001F807C0000000038003C003800000000000000000000000000000000000;
             char00[13] <= 256'h000001F80780000000038003C003800000000000000000000000000000000000;
             char00[14] <= 256'h000001F00F80000000038003C003800000000000000000000000000000000000;
             char00[15] <= 256'h000000F00F000E0000038003C003800000000000000000000000000000000000;
             char00[16] <= 256'h000000601E001F0000038103C003800000000000000000000000000000000000;
             char00[17] <= 256'h000000001C003F8000038383C003800000000000000000000000000000000000;
             char00[18] <= 256'h03FFFFFFFFFFFFC01FFFFFC3C003800000000000000000000000000000000000;
             char00[19] <= 256'h01FFFFFFFFFFFFE00FFFFFE3C003800000000000000000000000000000000000;
             char00[20] <= 256'h00F80007C000000000078003C003800000000000000000000000000000000000;
             char00[21] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
             char00[22] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
             char00[23] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
             char00[24] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
             char00[25] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
             char00[26] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
             char00[27] <= 256'h00000007C0000000000FE003C003800000000000000000000000000000000000;
             char00[28] <= 256'h00000007C0000000001FBC03C003800000000000000000000000000000000000;
             char00[29] <= 256'h00000007C0000000001F9F03C003800000000000000000000000000000000000;
             char00[30] <= 256'h00000007C0000380001F8F83C003800000000000000000000000000000000000;
             char00[31] <= 256'h00000007C00007C0003F87C3C003800000000000000000000000000000000000;
             char00[32] <= 256'h00000007C0000FE0003B83E3C003800000000000000000000000000000000000;
             char00[33] <= 256'h1FFFFFFFFFFFFFF0003B81E3C003800000000000000000000000000000000000;
             char00[34] <= 256'h0FFFFFFFFFFFFFF8007B80E3C003800000000000000000000000000000000000;
             char00[35] <= 256'h07C0000FB8000000007380E3C003800000000000000000000000000000000000;
             char00[36] <= 256'h0000000FBC00000000738043C003800000000000000000000000000000000000;
             char00[37] <= 256'h0000001F9C00000000E38003C003800000000000000000000000000000000000;
             char00[38] <= 256'h0000001F1E00000000E38003C003800000000000000000000000000000000000;
             char00[39] <= 256'h0000001F1E00000001C380038003800000000000000000000000000000000000;
             char00[40] <= 256'h0000003F0F00000001C380038003800000000000000000000000000000000000;
             char00[41] <= 256'h0000003E0F000000038380038003800000000000000000000000000000000000;
             char00[42] <= 256'h0000007E07800000030380078003800000000000000000000000000000000000;
             char00[43] <= 256'h000000FC07C00000070380078003800000000000000000000000000000000000;
             char00[44] <= 256'h000000F803C00000060380070003806000000000000000000000000000000000;
             char00[45] <= 256'h000001F803E000000C0380070003806000000000000000000000000000000000;
             char00[46] <= 256'h000003F001F000000C03800F0003806000000000000000000000000000000000;
             char00[47] <= 256'h000007E000F800001803800E0003806000000000000000000000000000000000;
             char00[48] <= 256'h000007C000FC00001003800E0003806000000000000000000000000000000000;
             char00[49] <= 256'h00000F80007F00002003801C0003806000000000000000000000000000000000;
             char00[50] <= 256'h00003F00003F80000003801C0003806000000000000000000000000000000000;
             char00[51] <= 256'h00007E00001FE000000380380003806000000000000000000000000000000000;
             char00[52] <= 256'h0000FC00000FF000000380380003806000000000000000000000000000000000;
             char00[53] <= 256'h0001F8000007FC0000038070000380F000000000000000000000000000000000;
             char00[54] <= 256'h0007E0000003FF80000380E00003C0F800000000000000000000000000000000;
             char00[55] <= 256'h001FC0000001FFF0000380C00003FFF800000000000000000000000000000000;
             char00[56] <= 256'h003F00000000FFFC000381800003FFF000000000000000000000000000000000;
             char00[57] <= 256'h00FC000000003FF0000383000000FFE000000000000000000000000000000000;
             char00[58] <= 256'h03F0000000001FC0000386000000000000000000000000000000000000000000;
             char00[59] <= 256'h1F8000000000078000038C000000000000000000000000000000000000000000;
             char00[60] <= 256'h1E00000000000000000398000000000000000000000000000000000000000000;
             char00[61] <= 256'h0000000000000000000200000000000000000000000000000000000000000000;
             char00[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
             char00[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    3'b100: begin //�ֶ�
             char00[  0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
             char00[  1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
             char00[  2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
             char00[  3] <= 256'h0000000000000000000000000080000000000000000000000000000000000000;
             char00[  4] <= 256'h000000000001E0000000000000F0000000000000000000000000000000000000;
             char00[  5] <= 256'h000000000007F0000000000000F8000000000000000000000000000000000000;
             char00[  6] <= 256'h00000000007FF0000000000000F0000000000000000000000000000000000000;
             char00[  7] <= 256'h000000000FFFF8000000000000F0000000000000000000000000000000000000;
             char00[  8] <= 256'h00000003FFFFFC000000000000F0000000000000000000000000000000000000;
             char00[  9] <= 256'h000007FFFFFFFC000000006000F0000000000000000000000000000000000000;
             char00[10] <= 256'h007FFFFFFF800000000000F000F0000000000000000000000000000000000000;
             char00[11] <= 256'h01FFFFFFC000000007FFFFF800F0000000000000000000000000000000000000;
             char00[12] <= 256'h00E00007C000000003FFFFFC00F0000000000000000000000000000000000000;
             char00[13] <= 256'h00000007C00000000100000000F0000000000000000000000000000000000000;
             char00[14] <= 256'h00000007C00000000000000000F0000000000000000000000000000000000000;
             char00[15] <= 256'h00000007C00000000000000000F0000000000000000000000000000000000000;
             char00[16] <= 256'h00000007C00000000000000000F0000000000000000000000000000000000000;
             char00[17] <= 256'h00000007C00000000000000000F0018000000000000000000000000000000000;
             char00[18] <= 256'h00000007C000000000000001FFFFFFE000000000000000000000000000000000;
             char00[19] <= 256'h00000007C000E00000000000FFFFFFE000000000000000000000000000000000;
             char00[20] <= 256'h00000007C001F0000000000000F003C000000000000000000000000000000000;
             char00[21] <= 256'h00000007C003F8000000000000F0038000000000000000000000000000000000;
             char00[22] <= 256'h00FFFFFFFFFFFC000000000C00F0038000000000000000000000000000000000;
             char00[23] <= 256'h007FFFFFFFFFFE000000001E00F0038000000000000000000000000000000000;
             char00[24] <= 256'h003E0007C00000001FFFFFFF00F0038000000000000000000000000000000000;
             char00[25] <= 256'h00000007C00000000FFFFFFF80E0038000000000000000000000000000000000;
             char00[26] <= 256'h00000007C00000000001C00000E0038000000000000000000000000000000000;
             char00[27] <= 256'h00000007C00000000001E00000E0038000000000000000000000000000000000;
             char00[28] <= 256'h00000007C00000000001F00000E0038000000000000000000000000000000000;
             char00[29] <= 256'h00000007C00000000003F00000E0038000000000000000000000000000000000;
             char00[30] <= 256'h00000007C00000000003E00000E0038000000000000000000000000000000000;
             char00[31] <= 256'h00000007C00001800003C00000E0038000000000000000000000000000000000;
             char00[32] <= 256'h00000007C00003C00007800001E0038000000000000000000000000000000000;
             char00[33] <= 256'h00000007C00007E00007000001C0038000000000000000000000000000000000;
             char00[34] <= 256'h00000007C0000FF0000F000001C0038000000000000000000000000000000000;
             char00[35] <= 256'h3FFFFFFFFFFFFFF8000E020001C0038000000000000000000000000000000000;
             char00[36] <= 256'h1FFFFFFFFFFFFFFC001C030001C0038000000000000000000000000000000000;
             char00[37] <= 256'h0F800007C0000000001C018003C0038000000000000000000000000000000000;
             char00[38] <= 256'h00000007C0000000003800C00380038000000000000000000000000000000000;
             char00[39] <= 256'h00000007C0000000007000E00380038000000000000000000000000000000000;
             char00[40] <= 256'h00000007C0000000006000700780038000000000000000000000000000000000;
             char00[41] <= 256'h00000007C000000000E000780700038000000000000000000000000000000000;
             char00[42] <= 256'h00000007C000000000C0003C0700078000000000000000000000000000000000;
             char00[43] <= 256'h00000007C00000000180003E0E00078000000000000000000000000000000000;
             char00[44] <= 256'h00000007C0000000030003FE0E00078000000000000000000000000000000000;
             char00[45] <= 256'h00000007C00000000607FFDE1C00078000000000000000000000000000000000;
             char00[46] <= 256'h00000007C00000001FFFF81E1C00078000000000000000000000000000000000;
             char00[47] <= 256'h00000007C00000000FFF000E3800078000000000000000000000000000000000;
             char00[48] <= 256'h00000007C00000000FF0000E7800078000000000000000000000000000000000;
             char00[49] <= 256'h00000007C00000000780000C7000070000000000000000000000000000000000;
             char00[50] <= 256'h00000007C000000006000000E000070000000000000000000000000000000000;
             char00[51] <= 256'h00000007C000000000000001C000070000000000000000000000000000000000;
             char00[52] <= 256'h00000007C00000000000000380000F0000000000000000000000000000000000;
             char00[53] <= 256'h0000000FC00000000000000700400F0000000000000000000000000000000000;
             char00[54] <= 256'h00003FFFC00000000000000E007FFE0000000000000000000000000000000000;
             char00[55] <= 256'h00003FFFC00000000000001C001FFE0000000000000000000000000000000000;
             char00[56] <= 256'h000007FF80000000000000380007FC0000000000000000000000000000000000;
             char00[57] <= 256'h000001FF80000000000000600003FC0000000000000000000000000000000000;
             char00[58] <= 256'h0000007F00000000000000C00001F80000000000000000000000000000000000;
             char00[59] <= 256'h0000003E00000000000003000000E00000000000000000000000000000000000;
             char00[60] <= 256'h0000003C00000000000002000000800000000000000000000000000000000000;
             char00[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
             char00[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
             char00[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    3'b010: begin//���Զ�
           char00[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
           char00[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
           char00[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
           char00[3] <= 256'h0000000600000000000000080000000000000000008000000000000000000000;
           char00[4] <= 256'h00000007800000000000000F000000000000000000F000000000000000000000;
           char00[5] <= 256'h00000007E00000000000000FC00000000000000000F800000000000000000000;
           char00[6] <= 256'h00000007E00000000000001F800000000000000000F000000000000000000000;
           char00[7] <= 256'h00000007C00000000000001F000000000000000000F000000000000000000000;
           char00[8] <= 256'h00000007C00380000000001E000000000000000000F000000000000000000000;
           char00[9] <= 256'h00180007C003E0000000001C000000000000006000F000000000000000000000;
           char00[10] <= 256'h001E0007C007F0000000003800000000000000F000F000000000000000000000;
           char00[11] <= 256'h000F0007C007F800000000300000800007FFFFF800F000000000000000000000;
           char00[12] <= 256'h0007C007C00FF000000000700000C00003FFFFFC00F000000000000000000000;
           char00[13] <= 256'h0003E007C00FE000000600600001E0000100000000F000000000000000000000;
           char00[14] <= 256'h0003F807C01F80000007FFFFFFFFF8000000000000F000000000000000000000;
           char00[15] <= 256'h0001FC07C01F00000007FFFFFFFFF8000000000000F000000000000000000000;
           char00[16] <= 256'h0000FE07C03E0000000780000001E0000000000000F000000000000000000000;
           char00[17] <= 256'h00007E07C07C0000000780000001E0000000000000F001800000000000000000;
           char00[18] <= 256'h00007F07C0780000000780000001E00000000001FFFFFFE00000000000000000;
           char00[19] <= 256'h00003F07C0F00000000780000001E00000000000FFFFFFE00000000000000000;
           char00[20] <= 256'h00003F07C1E00000000780000001E0000000000000F003C00000000000000000;
           char00[21] <= 256'h00001E07C3C00000000780000001E0000000000000F003800000000000000000;
           char00[22] <= 256'h00001E07C3800000000780000001E0000000000C00F003800000000000000000;
           char00[23] <= 256'h00000C07C7001800000780000001E0000000001E00F003800000000000000000;
           char00[24] <= 256'h00000007C0003C00000780000001E0001FFFFFFF00F003800000000000000000;
           char00[25] <= 256'h00000007C0007E00000780000001E0000FFFFFFF80E003800000000000000000;
           char00[26] <= 256'h03FFFFFFFFFFFF00000780000001E0000001C00000E003800000000000000000;
           char00[27] <= 256'h01FFFFFFFFFFFF800007FFFFFFFFE0000001E00000E003800000000000000000;
           char00[28] <= 256'h00F80007C00000000007FFFFFFFFE0000001F00000E003800000000000000000;
           char00[29] <= 256'h00000007C0000000000780000001E0000003F00000E003800000000000000000;
           char00[30] <= 256'h00000007C0000000000780000001E0000003E00000E003800000000000000000;
           char00[31] <= 256'h00000007C0000000000780000001E0000003C00000E003800000000000000000;
           char00[32] <= 256'h00000007C0000000000780000001E0000007800001E003800000000000000000;
           char00[33] <= 256'h00000007C0000000000780000001E0000007000001C003800000000000000000;
           char00[34] <= 256'h00000007C0000000000780000001E000000F000001C003800000000000000000;
           char00[35] <= 256'h00000007C0000000000780000001E000000E020001C003800000000000000000;
           char00[36] <= 256'h00000007C0000380000780000001E000001C030001C003800000000000000000;
           char00[37] <= 256'h00000007C00007C0000780000001E000001C018003C003800000000000000000;
           char00[38] <= 256'h00000007C0000FE0000780000001E000003800C0038003800000000000000000;
           char00[39] <= 256'h1FFFFFFFFFFFFFF0000780000001E000007000E0038003800000000000000000;
           char00[40] <= 256'h0FFFFFFFFFFFFFF8000780000001E00000600070078003800000000000000000;
           char00[41] <= 256'h07C00007C00000000007FFFFFFFFE00000E00078070003800000000000000000;
           char00[42] <= 256'h00000007C00000000007FFFFFFFFE00000C0003C070007800000000000000000;
           char00[43] <= 256'h00000007C0000000000780000001E0000180003E0E0007800000000000000000;
           char00[44] <= 256'h00000007C0000000000780000001E000030003FE0E0007800000000000000000;
           char00[45] <= 256'h00000007C0000000000780000001E0000607FFDE1C0007800000000000000000;
           char00[46] <= 256'h00000007C0000000000780000001E0001FFFF81E1C0007800000000000000000;
           char00[47] <= 256'h00000007C0000000000780000001E0000FFF000E380007800000000000000000;
           char00[48] <= 256'h00000007C0000000000780000001E0000FF0000E780007800000000000000000;
           char00[49] <= 256'h00000007C0000000000780000001E0000780000C700007000000000000000000;
           char00[50] <= 256'h00000007C0000000000780000001E00006000000E00007000000000000000000;
           char00[51] <= 256'h00000007C0000000000780000001E00000000001C00007000000000000000000;
           char00[52] <= 256'h00000007C0000000000780000001E0000000000380000F000000000000000000;
           char00[53] <= 256'h00000007C0000000000780000001E0000000000700400F000000000000000000;
           char00[54] <= 256'h00000007C00000000007FFFFFFFFE0000000000E007FFE000000000000000000;
           char00[55] <= 256'h00000007C00000000007FFFFFFFFE0000000001C001FFE000000000000000000;
           char00[56] <= 256'h00000007C0000000000780000001E000000000380007FC000000000000000000;
           char00[57] <= 256'h00000007C0000000000780000001E000000000600003FC000000000000000000;
           char00[58] <= 256'h00000007C0000000000780000001E000000000C00001F8000000000000000000;
           char00[59] <= 256'h00000007C0000000000780000001E000000003000000E0000000000000000000;
           char00[60] <= 256'h0000000700000000000600000001000000000200000080000000000000000000;
           char00[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
           char00[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
           char00[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    3'b001: begin//ȫ�Զ�
            char00[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
            char00[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
            char00[2] <= 256'h0000000E00000000000000000000000000000000000000000000000000000000;
            char00[3] <= 256'h0000000F80000000000000080000000000000000008000000000000000000000;
            char00[4] <= 256'h0000001FC00000000000000F000000000000000000F000000000000000000000;
            char00[5] <= 256'h0000001FE00000000000000FC00000000000000000F800000000000000000000;
            char00[6] <= 256'h0000003F800000000000001F800000000000000000F000000000000000000000;
            char00[7] <= 256'h0000003FC00000000000001F000000000000000000F000000000000000000000;
            char00[8] <= 256'h0000007FC00000000000001E000000000000000000F000000000000000000000;
            char00[9] <= 256'h0000007EE00000000000001C000000000000006000F000000000000000000000;
            char00[10] <= 256'h000000FCF00000000000003800000000000000F000F000000000000000000000;
            char00[11] <= 256'h000001F878000000000000300000800007FFFFF800F000000000000000000000;
            char00[12] <= 256'h000001F83C000000000000700000C00003FFFFFC00F000000000000000000000;
            char00[13] <= 256'h000003F03E000000000600600001E0000100000000F000000000000000000000;
            char00[14] <= 256'h000007E01F0000000007FFFFFFFFF8000000000000F000000000000000000000;
            char00[15] <= 256'h000007C00F8000000007FFFFFFFFF8000000000000F000000000000000000000;
            char00[16] <= 256'h00000FC007C00000000780000001E0000000000000F000000000000000000000;
            char00[17] <= 256'h00001F8003E00000000780000001E0000000000000F001800000000000000000;
            char00[18] <= 256'h00003F0003F00000000780000001E00000000001FFFFFFE00000000000000000;
            char00[19] <= 256'h00003E0001FC0000000780000001E00000000000FFFFFFE00000000000000000;
            char00[20] <= 256'h00007C0000FE0000000780000001E0000000000000F003C00000000000000000;
            char00[21] <= 256'h0000F800007F8000000780000001E0000000000000F003800000000000000000;
            char00[22] <= 256'h0001F800003FE000000780000001E0000000000C00F003800000000000000000;
            char00[23] <= 256'h0003F000000FF800000780000001E0000000001E00F003800000000000000000;
            char00[24] <= 256'h0007C000000FFF00000780000001E0001FFFFFFF00F003800000000000000000;
            char00[25] <= 256'h000F8000003FFFF0000780000001E0000FFFFFFF80E003800000000000000000;
            char00[26] <= 256'h003FFFFFFFFFFFFC000780000001E0000001C00000E003800000000000000000;
            char00[27] <= 256'h007FFFFFFFFFFFF80007FFFFFFFFE0000001E00000E003800000000000000000;
            char00[28] <= 256'h00F9F007C0001FE00007FFFFFFFFE0000001F00000E003800000000000000000;
            char00[29] <= 256'h01F00007C0000780000780000001E0000003F00000E003800000000000000000;
            char00[30] <= 256'h07C00007C0000180000780000001E0000003E00000E003800000000000000000;
            char00[31] <= 256'h1F000007C0000000000780000001E0000003C00000E003800000000000000000;
            char00[32] <= 256'h3C000007C0000000000780000001E0000007800001E003800000000000000000;
            char00[33] <= 256'h30000007C0000000000780000001E0000007000001C003800000000000000000;
            char00[34] <= 256'h00000007C0000000000780000001E000000F000001C003800000000000000000;
            char00[35] <= 256'h00000007C0000000000780000001E000000E020001C003800000000000000000;
            char00[36] <= 256'h00000007C0000000000780000001E000001C030001C003800000000000000000;
            char00[37] <= 256'h00000007C0030000000780000001E000001C018003C003800000000000000000;
            char00[38] <= 256'h00000007C0078000000780000001E000003800C0038003800000000000000000;
            char00[39] <= 256'h00000007C00FC000000780000001E000007000E0038003800000000000000000;
            char00[40] <= 256'h000FFFFFFFFFE000000780000001E00000600070078003800000000000000000;
            char00[41] <= 256'h0007FFFFFFFFF0000007FFFFFFFFE00000E00078070003800000000000000000;
            char00[42] <= 256'h0003E007C00000000007FFFFFFFFE00000C0003C070007800000000000000000;
            char00[43] <= 256'h00000007C0000000000780000001E0000180003E0E0007800000000000000000;
            char00[44] <= 256'h00000007C0000000000780000001E000030003FE0E0007800000000000000000;
            char00[45] <= 256'h00000007C0000000000780000001E0000607FFDE1C0007800000000000000000;
            char00[46] <= 256'h00000007C0000000000780000001E0001FFFF81E1C0007800000000000000000;
            char00[47] <= 256'h00000007C0000000000780000001E0000FFF000E380007800000000000000000;
            char00[48] <= 256'h00000007C0000000000780000001E0000FF0000E780007800000000000000000;
            char00[49] <= 256'h00000007C0000000000780000001E0000780000C700007000000000000000000;
            char00[50] <= 256'h00000007C0000000000780000001E00006000000E00007000000000000000000;
            char00[51] <= 256'h00000007C0000000000780000001E00000000001C00007000000000000000000;
            char00[52] <= 256'h00000007C0000000000780000001E0000000000380000F000000000000000000;
            char00[53] <= 256'h00000007C0000700000780000001E0000000000700400F000000000000000000;
            char00[54] <= 256'h00000007C0000F800007FFFFFFFFE0000000000E007FFE000000000000000000;
            char00[55] <= 256'h00000007C0001FC00007FFFFFFFFE0000000001C001FFE000000000000000000;
            char00[56] <= 256'h0FFFFFFFFFFFFFE0000780000001E000000000380007FC000000000000000000;
            char00[57] <= 256'h07FFFFFFFFFFFFF0000780000001E000000000600003FC000000000000000000;
            char00[58] <= 256'h03E0000000000000000780000001E000000000C00001F8000000000000000000;
            char00[59] <= 256'h0000000000000000000780000001E000000003000000E0000000000000000000;
            char00[60] <= 256'h0000000000000000000600000001000000000200000080000000000000000000;
            char00[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
            char00[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
            char00[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    default: begin
                 char00[  0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
                 char00[  1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
                 char00[  2] <= 256'h0000000000000000000200000000000000000000000000000000000000000000;
                 char00[  3] <= 256'h0000600000E00000000380000000000000000000000000000000000000000000;
                 char00[  4] <= 256'h0000780000F800000003E0000000000000000000000000000000000000000000;
                 char00[  5] <= 256'h00003E0000FC00000003C0000000000000000000000000000000000000000000;
                 char00[  6] <= 256'h00001F0001FF0000000380000000000000000000000000000000000000000000;
                 char00[  7] <= 256'h00000F8001FE0000000380020001000000000000000000000000000000000000;
                 char00[  8] <= 256'h00000FC001F80000000380038003800000000000000000000000000000000000;
                 char00[  9] <= 256'h000007E003F0000000038003FFFFE00000000000000000000000000000000000;
                 char00[10] <= 256'h000003F003E0000000038003FFFFF00000000000000000000000000000000000;
                 char00[11] <= 256'h000003F803E0000000038003C003C00000000000000000000000000000000000;
                 char00[12] <= 256'h000001F807C0000000038003C003800000000000000000000000000000000000;
                 char00[13] <= 256'h000001F80780000000038003C003800000000000000000000000000000000000;
                 char00[14] <= 256'h000001F00F80000000038003C003800000000000000000000000000000000000;
                 char00[15] <= 256'h000000F00F000E0000038003C003800000000000000000000000000000000000;
                 char00[16] <= 256'h000000601E001F0000038103C003800000000000000000000000000000000000;
                 char00[17] <= 256'h000000001C003F8000038383C003800000000000000000000000000000000000;
                 char00[18] <= 256'h03FFFFFFFFFFFFC01FFFFFC3C003800000000000000000000000000000000000;
                 char00[19] <= 256'h01FFFFFFFFFFFFE00FFFFFE3C003800000000000000000000000000000000000;
                 char00[20] <= 256'h00F80007C000000000078003C003800000000000000000000000000000000000;
                 char00[21] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
                 char00[22] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
                 char00[23] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
                 char00[24] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
                 char00[25] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
                 char00[26] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
                 char00[27] <= 256'h00000007C0000000000FE003C003800000000000000000000000000000000000;
                 char00[28] <= 256'h00000007C0000000001FBC03C003800000000000000000000000000000000000;
                 char00[29] <= 256'h00000007C0000000001F9F03C003800000000000000000000000000000000000;
                 char00[30] <= 256'h00000007C0000380001F8F83C003800000000000000000000000000000000000;
                 char00[31] <= 256'h00000007C00007C0003F87C3C003800000000000000000000000000000000000;
                 char00[32] <= 256'h00000007C0000FE0003B83E3C003800000000000000000000000000000000000;
                 char00[33] <= 256'h1FFFFFFFFFFFFFF0003B81E3C003800000000000000000000000000000000000;
                 char00[34] <= 256'h0FFFFFFFFFFFFFF8007B80E3C003800000000000000000000000000000000000;
                 char00[35] <= 256'h07C0000FB8000000007380E3C003800000000000000000000000000000000000;
                 char00[36] <= 256'h0000000FBC00000000738043C003800000000000000000000000000000000000;
                 char00[37] <= 256'h0000001F9C00000000E38003C003800000000000000000000000000000000000;
                 char00[38] <= 256'h0000001F1E00000000E38003C003800000000000000000000000000000000000;
                 char00[39] <= 256'h0000001F1E00000001C380038003800000000000000000000000000000000000;
                 char00[40] <= 256'h0000003F0F00000001C380038003800000000000000000000000000000000000;
                 char00[41] <= 256'h0000003E0F000000038380038003800000000000000000000000000000000000;
                 char00[42] <= 256'h0000007E07800000030380078003800000000000000000000000000000000000;
                 char00[43] <= 256'h000000FC07C00000070380078003800000000000000000000000000000000000;
                 char00[44] <= 256'h000000F803C00000060380070003806000000000000000000000000000000000;
                 char00[45] <= 256'h000001F803E000000C0380070003806000000000000000000000000000000000;
                 char00[46] <= 256'h000003F001F000000C03800F0003806000000000000000000000000000000000;
                 char00[47] <= 256'h000007E000F800001803800E0003806000000000000000000000000000000000;
                 char00[48] <= 256'h000007C000FC00001003800E0003806000000000000000000000000000000000;
                 char00[49] <= 256'h00000F80007F00002003801C0003806000000000000000000000000000000000;
                 char00[50] <= 256'h00003F00003F80000003801C0003806000000000000000000000000000000000;
                 char00[51] <= 256'h00007E00001FE000000380380003806000000000000000000000000000000000;
                 char00[52] <= 256'h0000FC00000FF000000380380003806000000000000000000000000000000000;
                 char00[53] <= 256'h0001F8000007FC0000038070000380F000000000000000000000000000000000;
                 char00[54] <= 256'h0007E0000003FF80000380E00003C0F800000000000000000000000000000000;
                 char00[55] <= 256'h001FC0000001FFF0000380C00003FFF800000000000000000000000000000000;
                 char00[56] <= 256'h003F00000000FFFC000381800003FFF000000000000000000000000000000000;
                 char00[57] <= 256'h00FC000000003FF0000383000000FFE000000000000000000000000000000000;
                 char00[58] <= 256'h03F0000000001FC0000386000000000000000000000000000000000000000000;
                 char00[59] <= 256'h1F8000000000078000038C000000000000000000000000000000000000000000;
                 char00[60] <= 256'h1E00000000000000000398000000000000000000000000000000000000000000;
                 char00[61] <= 256'h0000000000000000000200000000000000000000000000000000000000000000;
                 char00[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
                 char00[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
 endcase
 
 case(state)
    off: begin//�ػ�
        char11[  0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[  1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[  2] <= 256'h0000000000000000000200000000000000000000000000000000000000000000;
        char11[  3] <= 256'h0000600000E00000000380000000000000000000000000000000000000000000;
        char11[  4] <= 256'h0000780000F800000003E0000000000000000000000000000000000000000000;
        char11[  5] <= 256'h00003E0000FC00000003C0000000000000000000000000000000000000000000;
        char11[  6] <= 256'h00001F0001FF0000000380000000000000000000000000000000000000000000;
        char11[  7] <= 256'h00000F8001FE0000000380020001000000000000000000000000000000000000;
        char11[  8] <= 256'h00000FC001F80000000380038003800000000000000000000000000000000000;
        char11[  9] <= 256'h000007E003F0000000038003FFFFE00000000000000000000000000000000000;
        char11[10] <= 256'h000003F003E0000000038003FFFFF00000000000000000000000000000000000;
        char11[11] <= 256'h000003F803E0000000038003C003C00000000000000000000000000000000000;
        char11[12] <= 256'h000001F807C0000000038003C003800000000000000000000000000000000000;
        char11[13] <= 256'h000001F80780000000038003C003800000000000000000000000000000000000;
        char11[14] <= 256'h000001F00F80000000038003C003800000000000000000000000000000000000;
        char11[15] <= 256'h000000F00F000E0000038003C003800000000000000000000000000000000000;
        char11[16] <= 256'h000000601E001F0000038103C003800000000000000000000000000000000000;
        char11[17] <= 256'h000000001C003F8000038383C003800000000000000000000000000000000000;
        char11[18] <= 256'h03FFFFFFFFFFFFC01FFFFFC3C003800000000000000000000000000000000000;
        char11[19] <= 256'h01FFFFFFFFFFFFE00FFFFFE3C003800000000000000000000000000000000000;
        char11[20] <= 256'h00F80007C000000000078003C003800000000000000000000000000000000000;
        char11[21] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
        char11[22] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
        char11[23] <= 256'h00000007C000000000078003C003800000000000000000000000000000000000;
        char11[24] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
        char11[25] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
        char11[26] <= 256'h00000007C0000000000F8003C003800000000000000000000000000000000000;
        char11[27] <= 256'h00000007C0000000000FE003C003800000000000000000000000000000000000;
        char11[28] <= 256'h00000007C0000000001FBC03C003800000000000000000000000000000000000;
        char11[29] <= 256'h00000007C0000000001F9F03C003800000000000000000000000000000000000;
        char11[30] <= 256'h00000007C0000380001F8F83C003800000000000000000000000000000000000;
        char11[31] <= 256'h00000007C00007C0003F87C3C003800000000000000000000000000000000000;
        char11[32] <= 256'h00000007C0000FE0003B83E3C003800000000000000000000000000000000000;
        char11[33] <= 256'h1FFFFFFFFFFFFFF0003B81E3C003800000000000000000000000000000000000;
        char11[34] <= 256'h0FFFFFFFFFFFFFF8007B80E3C003800000000000000000000000000000000000;
        char11[35] <= 256'h07C0000FB8000000007380E3C003800000000000000000000000000000000000;
        char11[36] <= 256'h0000000FBC00000000738043C003800000000000000000000000000000000000;
        char11[37] <= 256'h0000001F9C00000000E38003C003800000000000000000000000000000000000;
        char11[38] <= 256'h0000001F1E00000000E38003C003800000000000000000000000000000000000;
        char11[39] <= 256'h0000001F1E00000001C380038003800000000000000000000000000000000000;
        char11[40] <= 256'h0000003F0F00000001C380038003800000000000000000000000000000000000;
        char11[41] <= 256'h0000003E0F000000038380038003800000000000000000000000000000000000;
        char11[42] <= 256'h0000007E07800000030380078003800000000000000000000000000000000000;
        char11[43] <= 256'h000000FC07C00000070380078003800000000000000000000000000000000000;
        char11[44] <= 256'h000000F803C00000060380070003806000000000000000000000000000000000;
        char11[45] <= 256'h000001F803E000000C0380070003806000000000000000000000000000000000;
        char11[46] <= 256'h000003F001F000000C03800F0003806000000000000000000000000000000000;
        char11[47] <= 256'h000007E000F800001803800E0003806000000000000000000000000000000000;
        char11[48] <= 256'h000007C000FC00001003800E0003806000000000000000000000000000000000;
        char11[49] <= 256'h00000F80007F00002003801C0003806000000000000000000000000000000000;
        char11[50] <= 256'h00003F00003F80000003801C0003806000000000000000000000000000000000;
        char11[51] <= 256'h00007E00001FE000000380380003806000000000000000000000000000000000;
        char11[52] <= 256'h0000FC00000FF000000380380003806000000000000000000000000000000000;
        char11[53] <= 256'h0001F8000007FC0000038070000380F000000000000000000000000000000000;
        char11[54] <= 256'h0007E0000003FF80000380E00003C0F800000000000000000000000000000000;
        char11[55] <= 256'h001FC0000001FFF0000380C00003FFF800000000000000000000000000000000;
        char11[56] <= 256'h003F00000000FFFC000381800003FFF000000000000000000000000000000000;
        char11[57] <= 256'h00FC000000003FF0000383000000FFE000000000000000000000000000000000;
        char11[58] <= 256'h03F0000000001FC0000386000000000000000000000000000000000000000000;
        char11[59] <= 256'h1F8000000000078000038C000000000000000000000000000000000000000000;
        char11[60] <= 256'h1E00000000000000000398000000000000000000000000000000000000000000;
        char11[61] <= 256'h0000000000000000000200000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    no_st: begin//δ��
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0000000700000000000010000000000000000001000000000000000000000000;
        char11[3] <= 256'h00000007C000000000001C000000000000000001C00000000000000000000000;
        char11[4] <= 256'h00000007F000000000001F000000000000000001F80000000000000000000000;
        char11[5] <= 256'h00000007F800000000001E000000000000000001F00000000000000000000000;
        char11[6] <= 256'h00000007E000000000001C000000000000000001E00000000000000000000000;
        char11[7] <= 256'h00000007E000000000001C000000000000000001E00000000000000000000000;
        char11[8] <= 256'h00000007E000000000001C000000000000000001E00000000000000000000000;
        char11[9] <= 256'h00000007E000000000001C000000040000010001E00000000000000000000000;
        char11[10] <= 256'h00000007E000000000001C0400000F000001E001E00030000000000000000000;
        char11[11] <= 256'h00000007E001C00000001C0C1FFFFF800001F801E00078000000000000000000;
        char11[12] <= 256'h00000007E003E00000001C1E0FFFFF000001E001FFFFFC000000000000000000;
        char11[13] <= 256'h00000007E007F00001FFFFFF04000F000001E001FFFFFE000000000000000000;
        char11[14] <= 256'h003FFFFFFFFFF80000FFFFFF80000F000001E001E00000000000000000000000;
        char11[15] <= 256'h001FFFFFFFFFFC0000401C0000000F000001E001E00000000000000000000000;
        char11[16] <= 256'h000F8007E000000000001C0000000F000001E001E00000000000000000000000;
        char11[17] <= 256'h00000007E000000000001C0000000F000001E001E00000000000000000000000;
        char11[18] <= 256'h00000007E000000000001C0000000F000001E001E00000000000000000000000;
        char11[19] <= 256'h00000007E000000000001C0000000F000001E001E00000000000000000000000;
        char11[20] <= 256'h00000007E000000000001C0000000F000001E001E00000000000000000000000;
        char11[21] <= 256'h00000007E000000000001C0000000F000001E001E00000000000000000000000;
        char11[22] <= 256'h00000007E000000000001C0000000F000001E001E00001000000000000000000;
        char11[23] <= 256'h00000007E000000000001C0300000F000001E001E00003800000000000000000;
        char11[24] <= 256'h00000007E000000000001C078C000F000001E001E00007C00000000000000000;
        char11[25] <= 256'h00000007E0000F000FFFFFFFCFFFFF001FFFFFFFFFFFFFE00000000000000000;
        char11[26] <= 256'h00000007E0001F8007FFFFFFEFFFFF000FFFFFFFFFFFFFF00000000000000000;
        char11[27] <= 256'h00000007E0003FC002001C000F000F0006000002000000000000000000000000;
        char11[28] <= 256'h0FFFFFFFFFFFFFE000001F000F000F0000000001800000000000000000000000;
        char11[29] <= 256'h07FFFFFFFFFFFFF000001F000F000C0000000001E00000000000000000000000;
        char11[30] <= 256'h0380003FF800000000001E000F00000000000001F80000000000000000000000;
        char11[31] <= 256'h0000003FFC00000000001E000F00000000000001E00000000000000000000000;
        char11[32] <= 256'h0000007FFC00000000601E000F00000000002001E00000000000000000000000;
        char11[33] <= 256'h0000007FEE00000000781E000F00000000003001E00008000000000000000000;
        char11[34] <= 256'h000000FFEE000000007E1E000F0000C000003801E0001C000000000000000000;
        char11[35] <= 256'h000001FFEF000000007C1E000F0000C000007E01E0003E000000000000000000;
        char11[36] <= 256'h000001F7E780000000781E060F0000C00000FC01E0003F000000000000000000;
        char11[37] <= 256'h000003F7E780000000781E0F0F0000C00000F001E0007F000000000000000000;
        char11[38] <= 256'h000007E7E3C0000000781FFF8F0000C00001F001E000FC000000000000000000;
        char11[39] <= 256'h00000FC7E3E0000000781FFFCF0000C00001E001E001F8000000000000000000;
        char11[40] <= 256'h00001F87E1F0000000701E000F0000C00003C001E003F0000000000000000000;
        char11[41] <= 256'h00001F07E0F8000000701E000F0000C000078001E007E0000000000000000000;
        char11[42] <= 256'h00003E07E0FC000000701E000F0000C000070001E00FC0000000000000000000;
        char11[43] <= 256'h00007C07E07E000000F01E000F0000E0000F0001E01F00000000000000000000;
        char11[44] <= 256'h0000F807E03F800000F01E00070000E0001E0001E03E00000000000000000000;
        char11[45] <= 256'h0001F007E01FC00000F81E00070001F8001C0001E07C00000000000000000000;
        char11[46] <= 256'h0003E007E00FF00000E81E0007FFFFF000380001E1F800000000000000000000;
        char11[47] <= 256'h0007C007E007F80000EC1E0003FFFFE000700001E3E000000000000000000000;
        char11[48] <= 256'h001F8007E003FE0000C71E0001FFFFC000E0000107C000000000000000000000;
        char11[49] <= 256'h003E0007E001FFC001C39E000000000000C000001F8000000000000000000000;
        char11[50] <= 256'h007C0007E000FFF801C1DE0000000000018000003E0000000000000000000000;
        char11[51] <= 256'h00F80007E0007FFC0180FE000000000003000000FC0000000000000000000000;
        char11[52] <= 256'h03E00007E0003FE003807E000000000004000003F00000000000000000000000;
        char11[53] <= 256'h07800007E0000F8003003FC0000000000000000FC00000000000000000000000;
        char11[54] <= 256'h1E000007E000070003000FF8000000000000003F800000000000000000000000;
        char11[55] <= 256'h18000007E0000000060003FFF0000038000000FC000000000000000000000000;
        char11[56] <= 256'h00000007E0000000060000FFFFFFFFF0000007F0000000000000000000000000;
        char11[57] <= 256'h00000007E00000000C00001FFFFFFFC000003F80000000000000000000000000;
        char11[58] <= 256'h00000007E000000008000001FFFFFF800001F800000000000000000000000000;
        char11[59] <= 256'h00000007C00000001800000007FFFF80001F8000000000000000000000000000;
        char11[60] <= 256'h0000000700000000100000000000000003F80000000000000000000000000000;
        char11[61] <= 256'h000000000000000000000000000000000E000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    start: begin//��
          char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0000380000000000000000010000000000000000000000000000000000000000;
        char11[3] <= 256'h00003E000000000000000001C000000000000000000000000000000000000000;
        char11[4] <= 256'h00003F800000000000000001F800000000000000000000000000000000000000;
        char11[5] <= 256'h00003F000000000000000001F000000000000000000000000000000000000000;
        char11[6] <= 256'h00003E000000000000000001E000000000000000000000000000000000000000;
        char11[7] <= 256'h00003E000000000000000001E000000000000000000000000000000000000000;
        char11[8] <= 256'h00003E000000000000000001E000000000000000000000000000000000000000;
        char11[9] <= 256'h00003E0000000E0000010001E000000000000000000000000000000000000000;
        char11[10] <= 256'h00003E0400000F800001E001E000300000000000000000000000000000000000;
        char11[11] <= 256'h00003E0E3FFFFFC00001F801E000780000000000000000000000000000000000;
        char11[12] <= 256'h00003E3F1FFFFF800001E001FFFFFC0000000000000000000000000000000000;
        char11[13] <= 256'h03FFFFFF8F801F000001E001FFFFFE0000000000000000000000000000000000;
        char11[14] <= 256'h01FFFFFFC0001F000001E001E000000000000000000000000000000000000000;
        char11[15] <= 256'h00F03E0000001F000001E001E000000000000000000000000000000000000000;
        char11[16] <= 256'h00003E0000001F000001E001E000000000000000000000000000000000000000;
        char11[17] <= 256'h00003E0000001F000001E001E000000000000000000000000000000000000000;
        char11[18] <= 256'h00003E0000001F000001E001E000000000000000000000000000000000000000;
        char11[19] <= 256'h00003E0000001F000001E001E000000000000000000000000000000000000000;
        char11[20] <= 256'h00003E0000001F000001E001E000000000000000000000000000000000000000;
        char11[21] <= 256'h00003E0000001F000001E001E000000000000000000000000000000000000000;
        char11[22] <= 256'h00003E0300001F000001E001E000010000000000000000000000000000000000;
        char11[23] <= 256'h00003E0788001F000001E001E000038000000000000000000000000000000000;
        char11[24] <= 256'h00003E0FCE001F000001E001E00007C000000000000000000000000000000000;
        char11[25] <= 256'h1FFFFFFFEFFFFF001FFFFFFFFFFFFFE000000000000000000000000000000000;
        char11[26] <= 256'h0FFFFFFFFFFFFF000FFFFFFFFFFFFFF000000000000000000000000000000000;
        char11[27] <= 256'h07801E000F801F00060000020000000000000000000000000000000000000000;
        char11[28] <= 256'h00001F800F801F00000000018000000000000000000000000000000000000000;
        char11[29] <= 256'h00001F800F801E0000000001E000000000000000000000000000000000000000;
        char11[30] <= 256'h00001F000F80000000000001F800000000000000000000000000000000000000;
        char11[31] <= 256'h00001F000F80000000000001E000000000000000000000000000000000000000;
        char11[32] <= 256'h00701F000F80000000002001E000000000000000000000000000000000000000;
        char11[33] <= 256'h007C1F000F80000000003001E000080000000000000000000000000000000000;
        char11[34] <= 256'h007F1F000F8000E000003801E0001C0000000000000000000000000000000000;
        char11[35] <= 256'h007E1F060F8000E000007E01E0003E0000000000000000000000000000000000;
        char11[36] <= 256'h00FC1F0F0F8000E00000FC01E0003F0000000000000000000000000000000000;
        char11[37] <= 256'h00FC1F1F8F8000E00000F001E0007F0000000000000000000000000000000000;
        char11[38] <= 256'h00FC1FFFCF8000E00001F001E000FC0000000000000000000000000000000000;
        char11[39] <= 256'h00F81FFFEF8000E00001E001E001F80000000000000000000000000000000000;
        char11[40] <= 256'h00F81F000F8000E00003C001E003F00000000000000000000000000000000000;
        char11[41] <= 256'h00F81F000F8001E000078001E007E00000000000000000000000000000000000;
        char11[42] <= 256'h00F81F000F0001E000070001E00FC00000000000000000000000000000000000;
        char11[43] <= 256'h00F81F000F0001F0000F0001E01F000000000000000000000000000000000000;
        char11[44] <= 256'h00F81F000F8001F0001E0001E03E000000000000000000000000000000000000;
        char11[45] <= 256'h01F81F000F8003FC001C0001E07C000000000000000000000000000000000000;
        char11[46] <= 256'h01FC1F000FFFFFF800380001E1F8000000000000000000000000000000000000;
        char11[47] <= 256'h01FE1F0007FFFFF000700001E3E0000000000000000000000000000000000000;
        char11[48] <= 256'h01EF1F0003FFFFE000E0000107C0000000000000000000000000000000000000;
        char11[49] <= 256'h01E7DF000000000000C000001F80000000000000000000000000000000000000;
        char11[50] <= 256'h03C3FF0000000000018000003E00000000000000000000000000000000000000;
        char11[51] <= 256'h03C1FF000000000003000000FC00000000000000000000000000000000000000;
        char11[52] <= 256'h03C0FF000000000004000003F000000000000000000000000000000000000000;
        char11[53] <= 256'h07807FE0000000000000000FC000000000000000000000000000000000000000;
        char11[54] <= 256'h07801FFF000000000000003F8000000000000000000000000000000000000000;
        char11[55] <= 256'h0F0007FFFFF03FFC000000FC0000000000000000000000000000000000000000;
        char11[56] <= 256'h0E0001FFFFFFFFF8000007F00000000000000000000000000000000000000000;
        char11[57] <= 256'h0E00003FFFFFFFE000003F800000000000000000000000000000000000000000;
        char11[58] <= 256'h1C000007FFFFFFC00001F8000000000000000000000000000000000000000000;
        char11[59] <= 256'h180000003FFFFF80001F80000000000000000000000000000000000000000000;
        char11[60] <= 256'h380000000007FF8003F800000000000000000000000000000000000000000000;
        char11[61] <= 256'h00000000000000000E0000000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    movef: begin//�ƶ�
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[3] <= 256'h0000000001C00000000000000080000000000000000000000000000000000000;
        char11[4] <= 256'h0000018001E000000000000000F0000000000000000000000000000000000000;
        char11[5] <= 256'h000007C003F000000000000000F8000000000000000000000000000000000000;
        char11[6] <= 256'h00001FE003F800000000000000F0000000000000000000000000000000000000;
        char11[7] <= 256'h0000FFE007E000000000000000F0000000000000000000000000000000000000;
        char11[8] <= 256'h0007FFF007C000000000000000F0000000000000000000000000000000000000;
        char11[9] <= 256'h007FFF000F8006000000006000F0000000000000000000000000000000000000;
        char11[10] <= 256'h07FFF0001F000F00000000F000F0000000000000000000000000000000000000;
        char11[11] <= 256'h0FF1F0001FFFFF8007FFFFF800F0000000000000000000000000000000000000;
        char11[12] <= 256'h0001F0003FFFFFC003FFFFFC00F0000000000000000000000000000000000000;
        char11[13] <= 256'h0001F0003C001FC00100000000F0000000000000000000000000000000000000;
        char11[14] <= 256'h0001F00078003F000000000000F0000000000000000000000000000000000000;
        char11[15] <= 256'h0001F000FE003E000000000000F0000000000000000000000000000000000000;
        char11[16] <= 256'h0001F001EF807C000000000000F0000000000000000000000000000000000000;
        char11[17] <= 256'h0001F003C7C0F8000000000000F0018000000000000000000000000000000000;
        char11[18] <= 256'h0001F00787E1F80000000001FFFFFFE000000000000000000000000000000000;
        char11[19] <= 256'h0001F00F03E3F00000000000FFFFFFE000000000000000000000000000000000;
        char11[20] <= 256'h0001F0EE03E7E0000000000000F003C000000000000000000000000000000000;
        char11[21] <= 256'h0001F1F003EFC0000000000000F0038000000000000000000000000000000000;
        char11[22] <= 256'h3FFFFFF801DF80000000000C00F0038000000000000000000000000000000000;
        char11[23] <= 256'h1FFFFFFC003F00000000001E00F0038000000000000000000000000000000000;
        char11[24] <= 256'h0F83F000007E00001FFFFFFF00F0038000000000000000000000000000000000;
        char11[25] <= 256'h0003F00001F800000FFFFFFF80E0038000000000000000000000000000000000;
        char11[26] <= 256'h0003F00003F000000001C00000E0038000000000000000000000000000000000;
        char11[27] <= 256'h0007F00007EE00000001E00000E0038000000000000000000000000000000000;
        char11[28] <= 256'h0007F0000F9F00000001F00000E0038000000000000000000000000000000000;
        char11[29] <= 256'h000FF0003F1F80000003F00000E0038000000000000000000000000000000000;
        char11[30] <= 256'h000FFC00FC3FC0000003E00000E0038000000000000000000000000000000000;
        char11[31] <= 256'h000FFF01F07F80000003C00000E0038000000000000000000000000000000000;
        char11[32] <= 256'h001FFF87C0FE00000007800001E0038000000000000000000000000000000000;
        char11[33] <= 256'h001FFFDF00FC00C00007000001C0038000000000000000000000000000000000;
        char11[34] <= 256'h003FF7FC01F801E0000F000001C0038000000000000000000000000000000000;
        char11[35] <= 256'h003FF3F003FFFFF0000E020001C0038000000000000000000000000000000000;
        char11[36] <= 256'h003FF3F007FFFFF8001C030001C0038000000000000000000000000000000000;
        char11[37] <= 256'h007FF1F00FC003F8001C018003C0038000000000000000000000000000000000;
        char11[38] <= 256'h007BF1E01F8007E0003800C00380038000000000000000000000000000000000;
        char11[39] <= 256'h00F3F0E03F000FC0007000E00380038000000000000000000000000000000000;
        char11[40] <= 256'h00F3F0007C000FC0006000700780038000000000000000000000000000000000;
        char11[41] <= 256'h01E3F000FE001F8000E000780700038000000000000000000000000000000000;
        char11[42] <= 256'h01C3F001FF803F0000C0003C0700078000000000000000000000000000000000;
        char11[43] <= 256'h03C3F007C7C03E000180003E0E00078000000000000000000000000000000000;
        char11[44] <= 256'h0783F00F87C07C00030003FE0E00078000000000000000000000000000000000;
        char11[45] <= 256'h0703F01E03E0FC000607FFDE1C00078000000000000000000000000000000000;
        char11[46] <= 256'h0E03F07C03E1F8001FFFF81E1C00078000000000000000000000000000000000;
        char11[47] <= 256'h0E03F07003E3F0000FFF000E3800078000000000000000000000000000000000;
        char11[48] <= 256'h1C03F00001E7E0000FF0000E7800078000000000000000000000000000000000;
        char11[49] <= 256'h3803F00001CFC0000780000C7000070000000000000000000000000000000000;
        char11[50] <= 256'h0003F000003F800006000000E000070000000000000000000000000000000000;
        char11[51] <= 256'h0003F000007F000000000001C000070000000000000000000000000000000000;
        char11[52] <= 256'h0003F00001FC00000000000380000F0000000000000000000000000000000000;
        char11[53] <= 256'h0003F00007F800000000000700400F0000000000000000000000000000000000;
        char11[54] <= 256'h0003F0000FE000000000000E007FFE0000000000000000000000000000000000;
        char11[55] <= 256'h0003F0007F8000000000001C001FFE0000000000000000000000000000000000;
        char11[56] <= 256'h0003F001FE000000000000380007FC0000000000000000000000000000000000;
        char11[57] <= 256'h0003F00FF8000000000000600003FC0000000000000000000000000000000000;
        char11[58] <= 256'h0003F07FC0000000000000C00001F80000000000000000000000000000000000;
        char11[59] <= 256'h0003E7FC00000000000003000000E00000000000000000000000000000000000;
        char11[60] <= 256'h00038F8000000000000002000000800000000000000000000000000000000000;
        char11[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    moveb: begin
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[3] <= 256'h0000000001C00000000000000080000000000000000000000000000000000000;
        char11[4] <= 256'h0000018001E000000000000000F0000000000000000000000000000000000000;
        char11[5] <= 256'h000007C003F000000000000000F8000000000000000000000000000000000000;
        char11[6] <= 256'h00001FE003F800000000000000F0000000000000000000000000000000000000;
        char11[7] <= 256'h0000FFE007E000000000000000F0000000000000000000000000000000000000;
        char11[8] <= 256'h0007FFF007C000000000000000F0000000000000000000000000000000000000;
        char11[9] <= 256'h007FFF000F8006000000006000F0000000000000000000000000000000000000;
        char11[10] <= 256'h07FFF0001F000F00000000F000F0000000000000000000000000000000000000;
        char11[11] <= 256'h0FF1F0001FFFFF8007FFFFF800F0000000000000000000000000000000000000;
        char11[12] <= 256'h0001F0003FFFFFC003FFFFFC00F0000000000000000000000000000000000000;
        char11[13] <= 256'h0001F0003C001FC00100000000F0000000000000000000000000000000000000;
        char11[14] <= 256'h0001F00078003F000000000000F0000000000000000000000000000000000000;
        char11[15] <= 256'h0001F000FE003E000000000000F0000000000000000000000000000000000000;
        char11[16] <= 256'h0001F001EF807C000000000000F0000000000000000000000000000000000000;
        char11[17] <= 256'h0001F003C7C0F8000000000000F0018000000000000000000000000000000000;
        char11[18] <= 256'h0001F00787E1F80000000001FFFFFFE000000000000000000000000000000000;
        char11[19] <= 256'h0001F00F03E3F00000000000FFFFFFE000000000000000000000000000000000;
        char11[20] <= 256'h0001F0EE03E7E0000000000000F003C000000000000000000000000000000000;
        char11[21] <= 256'h0001F1F003EFC0000000000000F0038000000000000000000000000000000000;
        char11[22] <= 256'h3FFFFFF801DF80000000000C00F0038000000000000000000000000000000000;
        char11[23] <= 256'h1FFFFFFC003F00000000001E00F0038000000000000000000000000000000000;
        char11[24] <= 256'h0F83F000007E00001FFFFFFF00F0038000000000000000000000000000000000;
        char11[25] <= 256'h0003F00001F800000FFFFFFF80E0038000000000000000000000000000000000;
        char11[26] <= 256'h0003F00003F000000001C00000E0038000000000000000000000000000000000;
        char11[27] <= 256'h0007F00007EE00000001E00000E0038000000000000000000000000000000000;
        char11[28] <= 256'h0007F0000F9F00000001F00000E0038000000000000000000000000000000000;
        char11[29] <= 256'h000FF0003F1F80000003F00000E0038000000000000000000000000000000000;
        char11[30] <= 256'h000FFC00FC3FC0000003E00000E0038000000000000000000000000000000000;
        char11[31] <= 256'h000FFF01F07F80000003C00000E0038000000000000000000000000000000000;
        char11[32] <= 256'h001FFF87C0FE00000007800001E0038000000000000000000000000000000000;
        char11[33] <= 256'h001FFFDF00FC00C00007000001C0038000000000000000000000000000000000;
        char11[34] <= 256'h003FF7FC01F801E0000F000001C0038000000000000000000000000000000000;
        char11[35] <= 256'h003FF3F003FFFFF0000E020001C0038000000000000000000000000000000000;
        char11[36] <= 256'h003FF3F007FFFFF8001C030001C0038000000000000000000000000000000000;
        char11[37] <= 256'h007FF1F00FC003F8001C018003C0038000000000000000000000000000000000;
        char11[38] <= 256'h007BF1E01F8007E0003800C00380038000000000000000000000000000000000;
        char11[39] <= 256'h00F3F0E03F000FC0007000E00380038000000000000000000000000000000000;
        char11[40] <= 256'h00F3F0007C000FC0006000700780038000000000000000000000000000000000;
        char11[41] <= 256'h01E3F000FE001F8000E000780700038000000000000000000000000000000000;
        char11[42] <= 256'h01C3F001FF803F0000C0003C0700078000000000000000000000000000000000;
        char11[43] <= 256'h03C3F007C7C03E000180003E0E00078000000000000000000000000000000000;
        char11[44] <= 256'h0783F00F87C07C00030003FE0E00078000000000000000000000000000000000;
        char11[45] <= 256'h0703F01E03E0FC000607FFDE1C00078000000000000000000000000000000000;
        char11[46] <= 256'h0E03F07C03E1F8001FFFF81E1C00078000000000000000000000000000000000;
        char11[47] <= 256'h0E03F07003E3F0000FFF000E3800078000000000000000000000000000000000;
        char11[48] <= 256'h1C03F00001E7E0000FF0000E7800078000000000000000000000000000000000;
        char11[49] <= 256'h3803F00001CFC0000780000C7000070000000000000000000000000000000000;
        char11[50] <= 256'h0003F000003F800006000000E000070000000000000000000000000000000000;
        char11[51] <= 256'h0003F000007F000000000001C000070000000000000000000000000000000000;
        char11[52] <= 256'h0003F00001FC00000000000380000F0000000000000000000000000000000000;
        char11[53] <= 256'h0003F00007F800000000000700400F0000000000000000000000000000000000;
        char11[54] <= 256'h0003F0000FE000000000000E007FFE0000000000000000000000000000000000;
        char11[55] <= 256'h0003F0007F8000000000001C001FFE0000000000000000000000000000000000;
        char11[56] <= 256'h0003F001FE000000000000380007FC0000000000000000000000000000000000;
        char11[57] <= 256'h0003F00FF8000000000000600003FC0000000000000000000000000000000000;
        char11[58] <= 256'h0003F07FC0000000000000C00001F80000000000000000000000000000000000;
        char11[59] <= 256'h0003E7FC00000000000003000000E00000000000000000000000000000000000;
        char11[60] <= 256'h00038F8000000000000002000000800000000000000000000000000000000000;
        char11[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;

    end
    semi_movef: begin
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[3] <= 256'h0000000001C00000000000000080000000000000000000000000000000000000;
        char11[4] <= 256'h0000018001E000000000000000F0000000000000000000000000000000000000;
        char11[5] <= 256'h000007C003F000000000000000F8000000000000000000000000000000000000;
        char11[6] <= 256'h00001FE003F800000000000000F0000000000000000000000000000000000000;
        char11[7] <= 256'h0000FFE007E000000000000000F0000000000000000000000000000000000000;
        char11[8] <= 256'h0007FFF007C000000000000000F0000000000000000000000000000000000000;
        char11[9] <= 256'h007FFF000F8006000000006000F0000000000000000000000000000000000000;
        char11[10] <= 256'h07FFF0001F000F00000000F000F0000000000000000000000000000000000000;
        char11[11] <= 256'h0FF1F0001FFFFF8007FFFFF800F0000000000000000000000000000000000000;
        char11[12] <= 256'h0001F0003FFFFFC003FFFFFC00F0000000000000000000000000000000000000;
        char11[13] <= 256'h0001F0003C001FC00100000000F0000000000000000000000000000000000000;
        char11[14] <= 256'h0001F00078003F000000000000F0000000000000000000000000000000000000;
        char11[15] <= 256'h0001F000FE003E000000000000F0000000000000000000000000000000000000;
        char11[16] <= 256'h0001F001EF807C000000000000F0000000000000000000000000000000000000;
        char11[17] <= 256'h0001F003C7C0F8000000000000F0018000000000000000000000000000000000;
        char11[18] <= 256'h0001F00787E1F80000000001FFFFFFE000000000000000000000000000000000;
        char11[19] <= 256'h0001F00F03E3F00000000000FFFFFFE000000000000000000000000000000000;
        char11[20] <= 256'h0001F0EE03E7E0000000000000F003C000000000000000000000000000000000;
        char11[21] <= 256'h0001F1F003EFC0000000000000F0038000000000000000000000000000000000;
        char11[22] <= 256'h3FFFFFF801DF80000000000C00F0038000000000000000000000000000000000;
        char11[23] <= 256'h1FFFFFFC003F00000000001E00F0038000000000000000000000000000000000;
        char11[24] <= 256'h0F83F000007E00001FFFFFFF00F0038000000000000000000000000000000000;
        char11[25] <= 256'h0003F00001F800000FFFFFFF80E0038000000000000000000000000000000000;
        char11[26] <= 256'h0003F00003F000000001C00000E0038000000000000000000000000000000000;
        char11[27] <= 256'h0007F00007EE00000001E00000E0038000000000000000000000000000000000;
        char11[28] <= 256'h0007F0000F9F00000001F00000E0038000000000000000000000000000000000;
        char11[29] <= 256'h000FF0003F1F80000003F00000E0038000000000000000000000000000000000;
        char11[30] <= 256'h000FFC00FC3FC0000003E00000E0038000000000000000000000000000000000;
        char11[31] <= 256'h000FFF01F07F80000003C00000E0038000000000000000000000000000000000;
        char11[32] <= 256'h001FFF87C0FE00000007800001E0038000000000000000000000000000000000;
        char11[33] <= 256'h001FFFDF00FC00C00007000001C0038000000000000000000000000000000000;
        char11[34] <= 256'h003FF7FC01F801E0000F000001C0038000000000000000000000000000000000;
        char11[35] <= 256'h003FF3F003FFFFF0000E020001C0038000000000000000000000000000000000;
        char11[36] <= 256'h003FF3F007FFFFF8001C030001C0038000000000000000000000000000000000;
        char11[37] <= 256'h007FF1F00FC003F8001C018003C0038000000000000000000000000000000000;
        char11[38] <= 256'h007BF1E01F8007E0003800C00380038000000000000000000000000000000000;
        char11[39] <= 256'h00F3F0E03F000FC0007000E00380038000000000000000000000000000000000;
        char11[40] <= 256'h00F3F0007C000FC0006000700780038000000000000000000000000000000000;
        char11[41] <= 256'h01E3F000FE001F8000E000780700038000000000000000000000000000000000;
        char11[42] <= 256'h01C3F001FF803F0000C0003C0700078000000000000000000000000000000000;
        char11[43] <= 256'h03C3F007C7C03E000180003E0E00078000000000000000000000000000000000;
        char11[44] <= 256'h0783F00F87C07C00030003FE0E00078000000000000000000000000000000000;
        char11[45] <= 256'h0703F01E03E0FC000607FFDE1C00078000000000000000000000000000000000;
        char11[46] <= 256'h0E03F07C03E1F8001FFFF81E1C00078000000000000000000000000000000000;
        char11[47] <= 256'h0E03F07003E3F0000FFF000E3800078000000000000000000000000000000000;
        char11[48] <= 256'h1C03F00001E7E0000FF0000E7800078000000000000000000000000000000000;
        char11[49] <= 256'h3803F00001CFC0000780000C7000070000000000000000000000000000000000;
        char11[50] <= 256'h0003F000003F800006000000E000070000000000000000000000000000000000;
        char11[51] <= 256'h0003F000007F000000000001C000070000000000000000000000000000000000;
        char11[52] <= 256'h0003F00001FC00000000000380000F0000000000000000000000000000000000;
        char11[53] <= 256'h0003F00007F800000000000700400F0000000000000000000000000000000000;
        char11[54] <= 256'h0003F0000FE000000000000E007FFE0000000000000000000000000000000000;
        char11[55] <= 256'h0003F0007F8000000000001C001FFE0000000000000000000000000000000000;
        char11[56] <= 256'h0003F001FE000000000000380007FC0000000000000000000000000000000000;
        char11[57] <= 256'h0003F00FF8000000000000600003FC0000000000000000000000000000000000;
        char11[58] <= 256'h0003F07FC0000000000000C00001F80000000000000000000000000000000000;
        char11[59] <= 256'h0003E7FC00000000000003000000E00000000000000000000000000000000000;
        char11[60] <= 256'h00038F8000000000000002000000800000000000000000000000000000000000;
        char11[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    keep_go: begin
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[3] <= 256'h0000000001C00000000000000080000000000000000000000000000000000000;
        char11[4] <= 256'h0000018001E000000000000000F0000000000000000000000000000000000000;
        char11[5] <= 256'h000007C003F000000000000000F8000000000000000000000000000000000000;
        char11[6] <= 256'h00001FE003F800000000000000F0000000000000000000000000000000000000;
        char11[7] <= 256'h0000FFE007E000000000000000F0000000000000000000000000000000000000;
        char11[8] <= 256'h0007FFF007C000000000000000F0000000000000000000000000000000000000;
        char11[9] <= 256'h007FFF000F8006000000006000F0000000000000000000000000000000000000;
        char11[10] <= 256'h07FFF0001F000F00000000F000F0000000000000000000000000000000000000;
        char11[11] <= 256'h0FF1F0001FFFFF8007FFFFF800F0000000000000000000000000000000000000;
        char11[12] <= 256'h0001F0003FFFFFC003FFFFFC00F0000000000000000000000000000000000000;
        char11[13] <= 256'h0001F0003C001FC00100000000F0000000000000000000000000000000000000;
        char11[14] <= 256'h0001F00078003F000000000000F0000000000000000000000000000000000000;
        char11[15] <= 256'h0001F000FE003E000000000000F0000000000000000000000000000000000000;
        char11[16] <= 256'h0001F001EF807C000000000000F0000000000000000000000000000000000000;
        char11[17] <= 256'h0001F003C7C0F8000000000000F0018000000000000000000000000000000000;
        char11[18] <= 256'h0001F00787E1F80000000001FFFFFFE000000000000000000000000000000000;
        char11[19] <= 256'h0001F00F03E3F00000000000FFFFFFE000000000000000000000000000000000;
        char11[20] <= 256'h0001F0EE03E7E0000000000000F003C000000000000000000000000000000000;
        char11[21] <= 256'h0001F1F003EFC0000000000000F0038000000000000000000000000000000000;
        char11[22] <= 256'h3FFFFFF801DF80000000000C00F0038000000000000000000000000000000000;
        char11[23] <= 256'h1FFFFFFC003F00000000001E00F0038000000000000000000000000000000000;
        char11[24] <= 256'h0F83F000007E00001FFFFFFF00F0038000000000000000000000000000000000;
        char11[25] <= 256'h0003F00001F800000FFFFFFF80E0038000000000000000000000000000000000;
        char11[26] <= 256'h0003F00003F000000001C00000E0038000000000000000000000000000000000;
        char11[27] <= 256'h0007F00007EE00000001E00000E0038000000000000000000000000000000000;
        char11[28] <= 256'h0007F0000F9F00000001F00000E0038000000000000000000000000000000000;
        char11[29] <= 256'h000FF0003F1F80000003F00000E0038000000000000000000000000000000000;
        char11[30] <= 256'h000FFC00FC3FC0000003E00000E0038000000000000000000000000000000000;
        char11[31] <= 256'h000FFF01F07F80000003C00000E0038000000000000000000000000000000000;
        char11[32] <= 256'h001FFF87C0FE00000007800001E0038000000000000000000000000000000000;
        char11[33] <= 256'h001FFFDF00FC00C00007000001C0038000000000000000000000000000000000;
        char11[34] <= 256'h003FF7FC01F801E0000F000001C0038000000000000000000000000000000000;
        char11[35] <= 256'h003FF3F003FFFFF0000E020001C0038000000000000000000000000000000000;
        char11[36] <= 256'h003FF3F007FFFFF8001C030001C0038000000000000000000000000000000000;
        char11[37] <= 256'h007FF1F00FC003F8001C018003C0038000000000000000000000000000000000;
        char11[38] <= 256'h007BF1E01F8007E0003800C00380038000000000000000000000000000000000;
        char11[39] <= 256'h00F3F0E03F000FC0007000E00380038000000000000000000000000000000000;
        char11[40] <= 256'h00F3F0007C000FC0006000700780038000000000000000000000000000000000;
        char11[41] <= 256'h01E3F000FE001F8000E000780700038000000000000000000000000000000000;
        char11[42] <= 256'h01C3F001FF803F0000C0003C0700078000000000000000000000000000000000;
        char11[43] <= 256'h03C3F007C7C03E000180003E0E00078000000000000000000000000000000000;
        char11[44] <= 256'h0783F00F87C07C00030003FE0E00078000000000000000000000000000000000;
        char11[45] <= 256'h0703F01E03E0FC000607FFDE1C00078000000000000000000000000000000000;
        char11[46] <= 256'h0E03F07C03E1F8001FFFF81E1C00078000000000000000000000000000000000;
        char11[47] <= 256'h0E03F07003E3F0000FFF000E3800078000000000000000000000000000000000;
        char11[48] <= 256'h1C03F00001E7E0000FF0000E7800078000000000000000000000000000000000;
        char11[49] <= 256'h3803F00001CFC0000780000C7000070000000000000000000000000000000000;
        char11[50] <= 256'h0003F000003F800006000000E000070000000000000000000000000000000000;
        char11[51] <= 256'h0003F000007F000000000001C000070000000000000000000000000000000000;
        char11[52] <= 256'h0003F00001FC00000000000380000F0000000000000000000000000000000000;
        char11[53] <= 256'h0003F00007F800000000000700400F0000000000000000000000000000000000;
        char11[54] <= 256'h0003F0000FE000000000000E007FFE0000000000000000000000000000000000;
        char11[55] <= 256'h0003F0007F8000000000001C001FFE0000000000000000000000000000000000;
        char11[56] <= 256'h0003F001FE000000000000380007FC0000000000000000000000000000000000;
        char11[57] <= 256'h0003F00FF8000000000000600003FC0000000000000000000000000000000000;
        char11[58] <= 256'h0003F07FC0000000000000C00001F80000000000000000000000000000000000;
        char11[59] <= 256'h0003E7FC00000000000003000000E00000000000000000000000000000000000;
        char11[60] <= 256'h00038F8000000000000002000000800000000000000000000000000000000000;
        char11[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;

    end
    wait_command: begin//�ȴ�ָ��
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0001800000C00000000000000400000000000000000000000000000200000000;
        char11[3] <= 256'h0003C00001F000000000E0000700000000020000000000000000000380000000;
        char11[4] <= 256'h0003F00001F800000000F00007E00000000380030000000000000007E0000000;
        char11[5] <= 256'h0003F80001FC00000000FC00078000000003E003C000000000000007E0000000;
        char11[6] <= 256'h0007F80003F800000001F000078000000003F003E000000000000007C0000000;
        char11[7] <= 256'h0007E00203F000000001E000078000000003C003C00010000000000FC0000000;
        char11[8] <= 256'h000FC00703E001C00003C000078000000003C003C00078000000000F60000000;
        char11[9] <= 256'h000FC00F87C003E00003C000078000000003C003C000FC000000001F30000000;
        char11[10] <= 256'h001FFFFFC7FFFFF000078000078030000003C003C001FE000000003E30000000;
        char11[11] <= 256'h001FFFFFEFFFFFF800070000078078000003C003C007FC000000003E18000000;
        char11[12] <= 256'h003F38000F0E0000000E00FFFFFFFC000003C003C01FC0000000007C1C000000;
        char11[13] <= 256'h003E3C001E0F0000001E007FFFFFFE000003C003C07F0000000000780C000000;
        char11[14] <= 256'h007C1E001E078000001C0000078000000003C003C1F80000000000F80E000000;
        char11[15] <= 256'h00F81F003C07C00000382000078000000003C183C7C00180000001F007000000;
        char11[16] <= 256'h00F01F807803E00000703800078000000003C3C3DE000180000001E003800000;
        char11[17] <= 256'h01E00F807003E00000E03C00078000001FFFFFE3F0000180000003E003800000;
        char11[18] <= 256'h03C00F83E003E00000C07E00078000000FFFFFF3C0000180000007C001C00000;
        char11[19] <= 256'h07800F83C003E00001807C00078000000603C003C00001800000078000E00000;
        char11[20] <= 256'h0F000F83F003E0000300F800078000000003C003C000018000000F0000F00000;
        char11[21] <= 256'h0E000703F801C0000600F000078000000003C003C000018000001E1800780000;
        char11[22] <= 256'h1C000003F00030000801F000078001800003C003C00001C000003C1C003E0000;
        char11[23] <= 256'h18000003F00078000001E000078003C00003C003C00003C00000780F001F0000;
        char11[24] <= 256'h00000003F000FC000003CFFFFFFFFFE00003C003C00003F00000F007800F8000;
        char11[25] <= 256'h001FFFFFFFFFFE00000387FFFFFFFFF00003C003FFFFFFE00001E003E007E000;
        char11[26] <= 256'h000FFFFFFFFFFF0000078200000000000003C021FFFFFFC00003C003F003F800;
        char11[27] <= 256'h0007C003F0000000000F8000000000000003C0C0FFFFFF8000078001F001FE00;
        char11[28] <= 256'h00000003F0000000000F8000000200000003C30000000000000E0000F800FF80;
        char11[29] <= 256'h00000003F0000000001F8000000380000003CE0000000000001C0000F8007FF8;
        char11[30] <= 256'h00000003F00000C0003F80000003E0000003FC00000000000078000078001FF8;
        char11[31] <= 256'h00000003F00001C0003F80000003C0000003F0000000000000E0000070000F80;
        char11[32] <= 256'h00000003F00003E000778000000380000007E002000008000380000070020300;
        char11[33] <= 256'h1FFFFFFFFFFFFFF000E7800000038180001FC00300001E000600000000070000;
        char11[34] <= 256'h0FFFFFFFFFFFFFF800C78000000383C0007FC003FFFFFF001C000000000F8000;
        char11[35] <= 256'h07C0000000000000018783FFFFFFFFE001FFC003FFFFFF001007FFFFFFFFC000;
        char11[36] <= 256'h0000000000380000030781FFFFFFFFF007F3C003C0001E000003FFFFFFFFE000;
        char11[37] <= 256'h00000000003E000006078000000380000FE3C003C0001E0000010000001FC000;
        char11[38] <= 256'h00000000003F00000C078000000380000F83C003C0001E0000000000003F0000;
        char11[39] <= 256'h00000000003F818018078004000380000703C003C0001E0000000000003E0000;
        char11[40] <= 256'h00000000003E03C010078006000380000203C003C0001E000000000000780000;
        char11[41] <= 256'h00000000003E07E000078003800380000203C003C0001E000000000000F00000;
        char11[42] <= 256'h03FFFFFFFFFFFFF000078003C00380000003C003C0001E000000000000E00000;
        char11[43] <= 256'h01FFFFFFFFFFFFF800078001E00380000003C003C0001E000000000001C00000;
        char11[44] <= 256'h00F80000003E000000078000F00380000003C003FFFFFE000000000003800000;
        char11[45] <= 256'h00001C00003E000000078000F00380000003C003FFFFFE000000000003000000;
        char11[46] <= 256'h00000F00003E000000078000F80380000003C003C0001E000000180006000000;
        char11[47] <= 256'h00000F80003E000000078000780380000003C003C0001E0000000F000E000000;
        char11[48] <= 256'h000007C0003E000000078000700380000003C003C0001E00000003C01C000000;
        char11[49] <= 256'h000003E0003E000000078000700380000003C003C0001E00000000F818000000;
        char11[50] <= 256'h000003F0003E000000078000200380000003C003C0001E000000007E30000000;
        char11[51] <= 256'h000001F8003E000000078000000380000003C003C0001E000000001FE0000000;
        char11[52] <= 256'h000001F8003E000000078000000380000003C003C0001E000000000FE0000000;
        char11[53] <= 256'h000001F8003E000000078000000380000003C003C0001E0000000007F8000000;
        char11[54] <= 256'h000000F0003E000000078000000380000003C003FFFFFE0000000001FC000000;
        char11[55] <= 256'h000000F0703E0000000780000003800007FFC003FFFFFE0000000000FE000000;
        char11[56] <= 256'h00000000FFFE0000000780000FC7800000FFC003C0001E00000000007F000000;
        char11[57] <= 256'h000000001FFE00000007800003FF8000003F8003C0001E00000000003F000000;
        char11[58] <= 256'h0000000007FC00000007800000FF8000001F0003C0001E00000000001F800000;
        char11[59] <= 256'h0000000003FC000000078000003F0000000E000380001800000000000F800000;
        char11[60] <= 256'h0000000001F8000000060000001E000000040002000000000000000007000000;
        char11[61] <= 256'h0000000000F00000000000000008000000000000000000000000000003000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    left_turning: begin//ת��
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0006000000700000000000100000000000000000000000000000000000000000;
        char11[3] <= 256'h00078000007C00000000001C0000000000000000000000000000000000000000;
        char11[4] <= 256'h0007E000007E00000000001F0000000000000000000000000000000000000000;
        char11[5] <= 256'h000FE000007F00000000003F0000000000000000000000000000000000000000;
        char11[6] <= 256'h000FC000007E00000000003E0000000000000000000000000000000000000000;
        char11[7] <= 256'h000F8000007C00000000003C0000000000000000000000000000000000000000;
        char11[8] <= 256'h000F800000F80000000000380000000000000000000000000000000000000000;
        char11[9] <= 256'h000F800000F80000000000700000000000000000000000000000000000000000;
        char11[10] <= 256'h001F008000F80000000000700000000000000000000000000000000000000000;
        char11[11] <= 256'h001F01C000F80700000000600000000000000000000000000000000000000000;
        char11[12] <= 256'h001F03E001F00F00004000E00000040000000000000000000000000000000000;
        char11[13] <= 256'h3FFFFFF001F01F80006000C000000E0000000000000000000000000000000000;
        char11[14] <= 256'h1FFFFFFFFFFFFFC0007FFFFFFFFFFF8000000000000000000000000000000000;
        char11[15] <= 256'h0FBE0007FFFFFFE0007FFFFFFFFFFF8000000000000000000000000000000000;
        char11[16] <= 256'h003E0003E1F000000078000000000F0000000000000000000000000000000000;
        char11[17] <= 256'h003C000003E000000078000000000E0000000000000000000000000000000000;
        char11[18] <= 256'h007C000003E000000078000000000E0000000000000000000000000000000000;
        char11[19] <= 256'h007DC00003E000000078000000000E0000000000000000000000000000000000;
        char11[20] <= 256'h007DF80003E000000078000000000E0000000000000000000000000000000000;
        char11[21] <= 256'h00F9FC0007C000000078000000000E0000000000000000000000000000000000;
        char11[22] <= 256'h00F9F80007C000000078000000000E0000000000000000000000000000000000;
        char11[23] <= 256'h00F9F00007C000C00078000000000E0000000000000000000000000000000000;
        char11[24] <= 256'h01F1F00007C001E00078000000800E0000000000000000000000000000000000;
        char11[25] <= 256'h01F1F0000F8007F00078060001C00E0000000000000000000000000000000000;
        char11[26] <= 256'h01F1F05FFFFFFFF8007807FFFFE00E0000000000000000000000000000000000;
        char11[27] <= 256'h03E1F0EFFFFFFFFC007807FFFFF00E0000000000000000000000000000000000;
        char11[28] <= 256'h07E1F1F7CF8000000078078001E00E0000000000000000000000000000000000;
        char11[29] <= 256'h0FFFFFF81F0000000078078001C00E0000000000000000000000000000000000;
        char11[30] <= 256'h07FFFFFC1F0000000078078001C00E0000000000000000000000000000000000;
        char11[31] <= 256'h03C1F0001F0000000078078001C00E0000000000000000000000000000000000;
        char11[32] <= 256'h0181F0003E0000000078078001C00E0000000000000000000000000000000000;
        char11[33] <= 256'h0001F0003E0000000078078001C00E0000000000000000000000000000000000;
        char11[34] <= 256'h0001F0007E0018000078078001C00E0000000000000000000000000000000000;
        char11[35] <= 256'h0001F0007C003C000078078001C00E0000000000000000000000000000000000;
        char11[36] <= 256'h0001F000FFFFFE000078078001C00E0000000000000000000000000000000000;
        char11[37] <= 256'h0001F000FFFFFF000078078001C00E0000000000000000000000000000000000;
        char11[38] <= 256'h0001F0067C007F800078078001C00E0000000000000000000000000000000000;
        char11[39] <= 256'h0001F0FE3800FF000078078001C00E0000000000000000000000000000000000;
        char11[40] <= 256'h0001FFF80000FC000078078001C00E0000000000000000000000000000000000;
        char11[41] <= 256'h0001FFC00001F800007807FFFFC00E0000000000000000000000000000000000;
        char11[42] <= 256'h001FFE000001F000007807FFFFC00E0000000000000000000000000000000000;
        char11[43] <= 256'h01FFF0000003E0000078078001C00E0000000000000000000000000000000000;
        char11[44] <= 256'h3FFFF0000003C0000078078001C00E0000000000000000000000000000000000;
        char11[45] <= 256'h3FFDF000000780000078078001C00E0000000000000000000000000000000000;
        char11[46] <= 256'h1FF1F000000780000078078001800E0000000000000000000000000000000000;
        char11[47] <= 256'h0F81F000F00F00000078060000000E0000000000000000000000000000000000;
        char11[48] <= 256'h0E01F0007E1E00000078000000000E0000000000000000000000000000000000;
        char11[49] <= 256'h0001F0001F9C00000078000000000E0000000000000000000000000000000000;
        char11[50] <= 256'h0001F0000FFC00000078000000000E0000000000000000000000000000000000;
        char11[51] <= 256'h0001F00003FC00000078000000000E0000000000000000000000000000000000;
        char11[52] <= 256'h0001F00001FF00000078000000000E0000000000000000000000000000000000;
        char11[53] <= 256'h0001F000007FC0000078000000001E0000000000000000000000000000000000;
        char11[54] <= 256'h0001F000003FE00000780000007FFE0000000000000000000000000000000000;
        char11[55] <= 256'h0001F000001FF00000780000001FFE0000000000000000000000000000000000;
        char11[56] <= 256'h0001F000000FF000007800000003FE0000000000000000000000000000000000;
        char11[57] <= 256'h0001F0000007F000007800000000FC0000000000000000000000000000000000;
        char11[58] <= 256'h0001F0000003F000007800000000780000000000000000000000000000000000;
        char11[59] <= 256'h0001F0000001F000007000000000700000000000000000000000000000000000;
        char11[60] <= 256'h0001E0000000E000004000000000000000000000000000000000000000000000;
        char11[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    right_turning: begin
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0006000000700000000000100000000000000000000000000000000000000000;
        char11[3] <= 256'h00078000007C00000000001C0000000000000000000000000000000000000000;
        char11[4] <= 256'h0007E000007E00000000001F0000000000000000000000000000000000000000;
        char11[5] <= 256'h000FE000007F00000000003F0000000000000000000000000000000000000000;
        char11[6] <= 256'h000FC000007E00000000003E0000000000000000000000000000000000000000;
        char11[7] <= 256'h000F8000007C00000000003C0000000000000000000000000000000000000000;
        char11[8] <= 256'h000F800000F80000000000380000000000000000000000000000000000000000;
        char11[9] <= 256'h000F800000F80000000000700000000000000000000000000000000000000000;
        char11[10] <= 256'h001F008000F80000000000700000000000000000000000000000000000000000;
        char11[11] <= 256'h001F01C000F80700000000600000000000000000000000000000000000000000;
        char11[12] <= 256'h001F03E001F00F00004000E00000040000000000000000000000000000000000;
        char11[13] <= 256'h3FFFFFF001F01F80006000C000000E0000000000000000000000000000000000;
        char11[14] <= 256'h1FFFFFFFFFFFFFC0007FFFFFFFFFFF8000000000000000000000000000000000;
        char11[15] <= 256'h0FBE0007FFFFFFE0007FFFFFFFFFFF8000000000000000000000000000000000;
        char11[16] <= 256'h003E0003E1F000000078000000000F0000000000000000000000000000000000;
        char11[17] <= 256'h003C000003E000000078000000000E0000000000000000000000000000000000;
        char11[18] <= 256'h007C000003E000000078000000000E0000000000000000000000000000000000;
        char11[19] <= 256'h007DC00003E000000078000000000E0000000000000000000000000000000000;
        char11[20] <= 256'h007DF80003E000000078000000000E0000000000000000000000000000000000;
        char11[21] <= 256'h00F9FC0007C000000078000000000E0000000000000000000000000000000000;
        char11[22] <= 256'h00F9F80007C000000078000000000E0000000000000000000000000000000000;
        char11[23] <= 256'h00F9F00007C000C00078000000000E0000000000000000000000000000000000;
        char11[24] <= 256'h01F1F00007C001E00078000000800E0000000000000000000000000000000000;
        char11[25] <= 256'h01F1F0000F8007F00078060001C00E0000000000000000000000000000000000;
        char11[26] <= 256'h01F1F05FFFFFFFF8007807FFFFE00E0000000000000000000000000000000000;
        char11[27] <= 256'h03E1F0EFFFFFFFFC007807FFFFF00E0000000000000000000000000000000000;
        char11[28] <= 256'h07E1F1F7CF8000000078078001E00E0000000000000000000000000000000000;
        char11[29] <= 256'h0FFFFFF81F0000000078078001C00E0000000000000000000000000000000000;
        char11[30] <= 256'h07FFFFFC1F0000000078078001C00E0000000000000000000000000000000000;
        char11[31] <= 256'h03C1F0001F0000000078078001C00E0000000000000000000000000000000000;
        char11[32] <= 256'h0181F0003E0000000078078001C00E0000000000000000000000000000000000;
        char11[33] <= 256'h0001F0003E0000000078078001C00E0000000000000000000000000000000000;
        char11[34] <= 256'h0001F0007E0018000078078001C00E0000000000000000000000000000000000;
        char11[35] <= 256'h0001F0007C003C000078078001C00E0000000000000000000000000000000000;
        char11[36] <= 256'h0001F000FFFFFE000078078001C00E0000000000000000000000000000000000;
        char11[37] <= 256'h0001F000FFFFFF000078078001C00E0000000000000000000000000000000000;
        char11[38] <= 256'h0001F0067C007F800078078001C00E0000000000000000000000000000000000;
        char11[39] <= 256'h0001F0FE3800FF000078078001C00E0000000000000000000000000000000000;
        char11[40] <= 256'h0001FFF80000FC000078078001C00E0000000000000000000000000000000000;
        char11[41] <= 256'h0001FFC00001F800007807FFFFC00E0000000000000000000000000000000000;
        char11[42] <= 256'h001FFE000001F000007807FFFFC00E0000000000000000000000000000000000;
        char11[43] <= 256'h01FFF0000003E0000078078001C00E0000000000000000000000000000000000;
        char11[44] <= 256'h3FFFF0000003C0000078078001C00E0000000000000000000000000000000000;
        char11[45] <= 256'h3FFDF000000780000078078001C00E0000000000000000000000000000000000;
        char11[46] <= 256'h1FF1F000000780000078078001800E0000000000000000000000000000000000;
        char11[47] <= 256'h0F81F000F00F00000078060000000E0000000000000000000000000000000000;
        char11[48] <= 256'h0E01F0007E1E00000078000000000E0000000000000000000000000000000000;
        char11[49] <= 256'h0001F0001F9C00000078000000000E0000000000000000000000000000000000;
        char11[50] <= 256'h0001F0000FFC00000078000000000E0000000000000000000000000000000000;
        char11[51] <= 256'h0001F00003FC00000078000000000E0000000000000000000000000000000000;
        char11[52] <= 256'h0001F00001FF00000078000000000E0000000000000000000000000000000000;
        char11[53] <= 256'h0001F000007FC0000078000000001E0000000000000000000000000000000000;
        char11[54] <= 256'h0001F000003FE00000780000007FFE0000000000000000000000000000000000;
        char11[55] <= 256'h0001F000001FF00000780000001FFE0000000000000000000000000000000000;
        char11[56] <= 256'h0001F000000FF000007800000003FE0000000000000000000000000000000000;
        char11[57] <= 256'h0001F0000007F000007800000000FC0000000000000000000000000000000000;
        char11[58] <= 256'h0001F0000003F000007800000000780000000000000000000000000000000000;
        char11[59] <= 256'h0001F0000001F000007000000000700000000000000000000000000000000000;
        char11[60] <= 256'h0001E0000000E000004000000000000000000000000000000000000000000000;
        char11[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;   
    end
    circle_turning: begin//��ͷ
        char11[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[3] <= 256'h0006000003800000000000004000000000000000000000000000000000000000;
        char11[4] <= 256'h0007800003E00000000000007000000000000000000000000000000000000000;
        char11[5] <= 256'h0007F00003F80000000000007C00000000000000000000000000000000000000;
        char11[6] <= 256'h0007E00003F80000000000007E00000000000000000000000000000000000000;
        char11[7] <= 256'h0007C00003F00000000000007C00000000000000000000000000000000000000;
        char11[8] <= 256'h0007C00003E000000001C0007800000000000000000000000000000000000000;
        char11[9] <= 256'h0007C00003E003800000F8007800000000000000000000000000000000000000;
        char11[10] <= 256'h0007C00003E007C000007E007800000000000000000000000000000000000000;
        char11[11] <= 256'h0007C00003FFFFE000003F807800000000000000000000000000000000000000;
        char11[12] <= 256'h0007C00003FFFFF000001FC07800000000000000000000000000000000000000;
        char11[13] <= 256'h0007C00003E0000000000FE07800000000000000000000000000000000000000;
        char11[14] <= 256'h0007C00003E00000000007E07800000000000000000000000000000000000000;
        char11[15] <= 256'h0007C30003E00000000003E07800000000000000000000000000000000000000;
        char11[16] <= 256'h0007C78003E00000000001E07800000000000000000000000000000000000000;
        char11[17] <= 256'h3FFFFFD803E00C00000001E07800000000000000000000000000000000000000;
        char11[18] <= 256'h1FFFFFFE03E01E00000000E07800000000000000000000000000000000000000;
        char11[19] <= 256'h0E07C01FFFFFFF00000000C07800000000000000000000000000000000000000;
        char11[20] <= 256'h0007C01FFFFFFF80007000007800000000000000000000000000000000000000;
        char11[21] <= 256'h0007C01F00003F00003C00007800000000000000000000000000000000000000;
        char11[22] <= 256'h0007C01F00003E00001F00007000000000000000000000000000000000000000;
        char11[23] <= 256'h0007C01F00003E00000FC0007000000000000000000000000000000000000000;
        char11[24] <= 256'h0007C01F00003E000007F0007000000000000000000000000000000000000000;
        char11[25] <= 256'h0007C01F00003E000003F0007000000000000000000000000000000000000000;
        char11[26] <= 256'h0007C05F00003E000001F8007000000000000000000000000000000000000000;
        char11[27] <= 256'h0007C1FF00003E000000F8007000000000000000000000000000000000000000;
        char11[28] <= 256'h0007CFDFFFFFFE000000F800F000000000000000000000000000000000000000;
        char11[29] <= 256'h0007FF1FFFFFFE0000007800F000000000000000000000000000000000000000;
        char11[30] <= 256'h0007FC1F00003E0000003800F000000000000000000000000000000000000000;
        char11[31] <= 256'h0007F81F00003E0000003000F000000000000000000000000000000000000000;
        char11[32] <= 256'h001FE01F00003E0000001000F000020000000000000000000000000000000000;
        char11[33] <= 256'h007FC01F00003E0000000000F000070000000000000000000000000000000000;
        char11[34] <= 256'h03FFC01F00003E0000000000F0000F8000000000000000000000000000000000;
        char11[35] <= 256'h1FFFC01F00003E0000000000F0001FC000000000000000000000000000000000;
        char11[36] <= 256'h1FF7C01F00003E000FFFFFFFFFFFFFE000000000000000000000000000000000;
        char11[37] <= 256'h1FC7C01FFFFFFE0007FFFFFFFFFFFFF000000000000000000000000000000000;
        char11[38] <= 256'h0F87C01FFFFFFE0002000001E000000000000000000000000000000000000000;
        char11[39] <= 256'h0607C01F03E03E0000000001E000000000000000000000000000000000000000;
        char11[40] <= 256'h0007C01F03E03E0000000001C000000000000000000000000000000000000000;
        char11[41] <= 256'h0007C01E03E0380000000003C000000000000000000000000000000000000000;
        char11[42] <= 256'h0007C01803E0000000000003C000000000000000000000000000000000000000;
        char11[43] <= 256'h0007C00003E0008000000007F000000000000000000000000000000000000000;
        char11[44] <= 256'h0007C00003E001C0000000079E00000000000000000000000000000000000000;
        char11[45] <= 256'h0007C00003E003E00000000F0F80000000000000000000000000000000000000;
        char11[46] <= 256'h0007DFFFFFFFFFF00000000F03E0000000000000000000000000000000000000;
        char11[47] <= 256'h0007CFFFFFFFFFF80000001E00FC000000000000000000000000000000000000;
        char11[48] <= 256'h0007C7C003E000000000003C007F000000000000000000000000000000000000;
        char11[49] <= 256'h0007C00003E0000000000078001FC00000000000000000000000000000000000;
        char11[50] <= 256'h0007C00003E00000000000F0000FF00000000000000000000000000000000000;
        char11[51] <= 256'h0007C00003E00000000001E00003FC0000000000000000000000000000000000;
        char11[52] <= 256'h0007C00003E00000000003C00001FE0000000000000000000000000000000000;
        char11[53] <= 256'h0007C00003E0000000000F8000007F8000000000000000000000000000000000;
        char11[54] <= 256'h0007C00003E0000000001F0000003F8000000000000000000000000000000000;
        char11[55] <= 256'h0FCFC00003E0000000007C0000001FC000000000000000000000000000000000;
        char11[56] <= 256'h07FF800003E000000001F00000000FC000000000000000000000000000000000;
        char11[57] <= 256'h01FF800003E000000007C000000007C000000000000000000000000000000000;
        char11[58] <= 256'h00FF800003E00000001E0000000003C000000000000000000000000000000000;
        char11[59] <= 256'h003F000003E0000000F80000000001C000000000000000000000000000000000;
        char11[60] <= 256'h001E000003E00000078000000000008000000000000000000000000000000000;
        char11[61] <= 256'h00180000038000000C0000000000000000000000000000000000000000000000;
        char11[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
        char11[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    end
    default: begin
        char11[0] <= char11[0];
        char11[1] <= char11[1];
        char11[2] <= char11[2];
        char11[3] <= char11[3];
        char11[4] <= char11[4];
        char11[5] <= char11[5];
        char11[6] <= char11[6];
        char11[7] <= char11[7];
        char11[8] <= char11[8];
        char11[9] <= char11[9];
        char11[10] <= char11[10];
        char11[11] <= char11[11];
        char11[12] <= char11[12];
        char11[13] <= char11[13];
        char11[14] <= char11[14];
        char11[15] <= char11[15];
        char11[16] <= char11[16];
        char11[17] <= char11[17];
        char11[18] <= char11[18];
        char11[19] <= char11[19];
        char11[20] <= char11[20];
        char11[21] <= char11[21];
        char11[22] <= char11[22];
        char11[23] <= char11[23];
        char11[24] <= char11[24];
        char11[25] <= char11[25];
        char11[26] <= char11[26];
        char11[27] <= char11[27];
        char11[28] <= char11[28];
        char11[29] <= char11[29];
        char11[30] <= char11[30];
        char11[31] <= char11[31];
        char11[32] <= char11[32];
        char11[33] <= char11[33];
        char11[34] <= char11[34];
        char11[35] <= char11[35];
        char11[36] <= char11[36];
        char11[37] <= char11[37];
        char11[38] <= char11[38];
        char11[39] <= char11[39];
        char11[40] <= char11[40];
        char11[41] <= char11[41];
        char11[42] <= char11[42];
        char11[43] <= char11[43];
        char11[44] <= char11[44];
        char11[45] <= char11[45];
        char11[46] <= char11[46];
        char11[47] <= char11[47];
        char11[48] <= char11[48];
        char11[49] <= char11[49];
        char11[50] <= char11[50];
        char11[51] <= char11[51];
        char11[52] <= char11[52];
        char11[53] <= char11[53];
        char11[54] <= char11[54];
        char11[55] <= char11[55];
        char11[56] <= char11[56];
        char11[57] <= char11[57];
        char11[58] <= char11[58];
        char11[59] <= char11[59];
        char11[60] <= char11[60];
        char11[61] <= char11[61];
        char11[62] <= char11[62];
        char11[63] <= char11[63];
    end
    
 endcase
 
 
         case(li/hkm)
             4'd0: begin
                 char22_0[  0] <= 32'h00000000;
                 char22_0[  1] <= 32'h00000000;
                 char22_0[  2] <= 32'h00000000;
                 char22_0[  3] <= 32'h00000000;
                 char22_0[  4] <= 32'h00000000;
                 char22_0[  5] <= 32'h00000000;
                 char22_0[  6] <= 32'h00000000;
                 char22_0[  7] <= 32'h00000000;
                 char22_0[  8] <= 32'h00000000;
                 char22_0[  9] <= 32'h00000000;
                 char22_0[10] <= 32'h000FF000;
                 char22_0[11] <= 32'h003FFC00;
                 char22_0[12] <= 32'h007E7E00;
                 char22_0[13] <= 32'h00F81F00;
                 char22_0[14] <= 32'h01F00F80;
                 char22_0[15] <= 32'h03F00FC0;
                 char22_0[16] <= 32'h03E007C0;
                 char22_0[17] <= 32'h07E007E0;
                 char22_0[18] <= 32'h07C003E0;
                 char22_0[19] <= 32'h0FC003F0;
                 char22_0[20] <= 32'h0FC003F0;
                 char22_0[21] <= 32'h0FC003F0;
                 char22_0[22] <= 32'h1F8001F8;
                 char22_0[23] <= 32'h1F8001F8;
                 char22_0[24] <= 32'h1F8001F8;
                 char22_0[25] <= 32'h1F8001F8;
                 char22_0[26] <= 32'h1F8001F8;
                 char22_0[27] <= 32'h3F8001F8;
                 char22_0[28] <= 32'h3F8001F8;
                 char22_0[29] <= 32'h3F8001F8;
                 char22_0[30] <= 32'h3F8001F8;
                 char22_0[31] <= 32'h3F8001F8;
                 char22_0[32] <= 32'h3F8001F8;
                 char22_0[33] <= 32'h3F8001F8;
                 char22_0[34] <= 32'h3F8001F8;
                 char22_0[35] <= 32'h3F8001F8;
                 char22_0[36] <= 32'h3F8001F8;
                 char22_0[37] <= 32'h1F8001F8;
                 char22_0[38] <= 32'h1F8001F8;
                 char22_0[39] <= 32'h1F8001F8;
                 char22_0[40] <= 32'h1F8001F8;
                 char22_0[41] <= 32'h1F8001F0;
                 char22_0[42] <= 32'h0F8003F0;
                 char22_0[43] <= 32'h0FC003F0;
                 char22_0[44] <= 32'h0FC003F0;
                 char22_0[45] <= 32'h07C003E0;
                 char22_0[46] <= 32'h07E007E0;
                 char22_0[47] <= 32'h03E007C0;
                 char22_0[48] <= 32'h03F00FC0;
                 char22_0[49] <= 32'h01F00F80;
                 char22_0[50] <= 32'h00F81F00;
                 char22_0[51] <= 32'h007E7E00;
                 char22_0[52] <= 32'h003FFC00;
                 char22_0[53] <= 32'h000FF000;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//0
             4'd1: begin
                 char22_0[  0] <= 32'h00000000;
                 char22_0[  1] <= 32'h00000000;
                 char22_0[  2] <= 32'h00000000;
                 char22_0[  3] <= 32'h00000000;
                 char22_0[  4] <= 32'h00000000;
                 char22_0[  5] <= 32'h00000000;
                 char22_0[  6] <= 32'h00000000;
                 char22_0[  7] <= 32'h00000000;
                 char22_0[  8] <= 32'h00000000;
                 char22_0[  9] <= 32'h00000000;
                 char22_0[10] <= 32'h0000E000;
                 char22_0[11] <= 32'h0001E000;
                 char22_0[12] <= 32'h0003E000;
                 char22_0[13] <= 32'h001FE000;
                 char22_0[14] <= 32'h03FFE000;
                 char22_0[15] <= 32'h03FFE000;
                 char22_0[16] <= 32'h0007E000;
                 char22_0[17] <= 32'h0007E000;
                 char22_0[18] <= 32'h0007E000;
                 char22_0[19] <= 32'h0007E000;
                 char22_0[20] <= 32'h0007E000;
                 char22_0[21] <= 32'h0007E000;
                 char22_0[22] <= 32'h0007E000;
                 char22_0[23] <= 32'h0007E000;
                 char22_0[24] <= 32'h0007E000;
                 char22_0[25] <= 32'h0007E000;
                 char22_0[26] <= 32'h0007E000;
                 char22_0[27] <= 32'h0007E000;
                 char22_0[28] <= 32'h0007E000;
                 char22_0[29] <= 32'h0007E000;
                 char22_0[30] <= 32'h0007E000;
                 char22_0[31] <= 32'h0007E000;
                 char22_0[32] <= 32'h0007E000;
                 char22_0[33] <= 32'h0007E000;
                 char22_0[34] <= 32'h0007E000;
                 char22_0[35] <= 32'h0007E000;
                 char22_0[36] <= 32'h0007E000;
                 char22_0[37] <= 32'h0007E000;
                 char22_0[38] <= 32'h0007E000;
                 char22_0[39] <= 32'h0007E000;
                 char22_0[40] <= 32'h0007E000;
                 char22_0[41] <= 32'h0007E000;
                 char22_0[42] <= 32'h0007E000;
                 char22_0[43] <= 32'h0007E000;
                 char22_0[44] <= 32'h0007E000;
                 char22_0[45] <= 32'h0007E000;
                 char22_0[46] <= 32'h0007E000;
                 char22_0[47] <= 32'h0007E000;
                 char22_0[48] <= 32'h0007E000;
                 char22_0[49] <= 32'h0007E000;
                 char22_0[50] <= 32'h0007E000;
                 char22_0[51] <= 32'h000FF800;
                 char22_0[52] <= 32'h03FFFFC0;
                 char22_0[53] <= 32'h03FFFFC0;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//1
             4'd2: begin
                 char22_0[  0] <= 32'h00000000;
                 char22_0[  1] <= 32'h00000000;
                 char22_0[  2] <= 32'h00000000;
                 char22_0[  3] <= 32'h00000000;
                 char22_0[  4] <= 32'h00000000;
                 char22_0[  5] <= 32'h00000000;
                 char22_0[  6] <= 32'h00000000;
                 char22_0[  7] <= 32'h00000000;
                 char22_0[  8] <= 32'h00000000;
                 char22_0[  9] <= 32'h00000000;
                 char22_0[10] <= 32'h001FFC00;
                 char22_0[11] <= 32'h007FFF00;
                 char22_0[12] <= 32'h01F83F80;
                 char22_0[13] <= 32'h03E00FC0;
                 char22_0[14] <= 32'h07C007E0;
                 char22_0[15] <= 32'h078007E0;
                 char22_0[16] <= 32'h0F8003F0;
                 char22_0[17] <= 32'h0F8003F0;
                 char22_0[18] <= 32'h1F8003F0;
                 char22_0[19] <= 32'h1F8003F0;
                 char22_0[20] <= 32'h1FC003F0;
                 char22_0[21] <= 32'h1FC003F0;
                 char22_0[22] <= 32'h1FC003F0;
                 char22_0[23] <= 32'h0FC003F0;
                 char22_0[24] <= 32'h07C003F0;
                 char22_0[25] <= 32'h000003E0;
                 char22_0[26] <= 32'h000007E0;
                 char22_0[27] <= 32'h000007E0;
                 char22_0[28] <= 32'h00000FC0;
                 char22_0[29] <= 32'h00000F80;
                 char22_0[30] <= 32'h00001F80;
                 char22_0[31] <= 32'h00003F00;
                 char22_0[32] <= 32'h00003E00;
                 char22_0[33] <= 32'h00007C00;
                 char22_0[34] <= 32'h0000F800;
                 char22_0[35] <= 32'h0001F000;
                 char22_0[36] <= 32'h0003E000;
                 char22_0[37] <= 32'h0007C000;
                 char22_0[38] <= 32'h000F8000;
                 char22_0[39] <= 32'h001F0000;
                 char22_0[40] <= 32'h003E0000;
                 char22_0[41] <= 32'h007C0000;
                 char22_0[42] <= 32'h00F80000;
                 char22_0[43] <= 32'h01F00038;
                 char22_0[44] <= 32'h01E00038;
                 char22_0[45] <= 32'h03C00070;
                 char22_0[46] <= 32'h07800070;
                 char22_0[47] <= 32'h0F8000F0;
                 char22_0[48] <= 32'h0F0000F0;
                 char22_0[49] <= 32'h1E0003F0;
                 char22_0[50] <= 32'h3FFFFFF0;
                 char22_0[51] <= 32'h3FFFFFF0;
                 char22_0[52] <= 32'h3FFFFFE0;
                 char22_0[53] <= 32'h3FFFFFE0;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//2
             4'd3: begin
                 char22_0[  0] <= 32'h00000000;
                 char22_0[  1] <= 32'h00000000;
                 char22_0[  2] <= 32'h00000000;
                 char22_0[  3] <= 32'h00000000;
                 char22_0[  4] <= 32'h00000000;
                 char22_0[  5] <= 32'h00000000;
                 char22_0[  6] <= 32'h00000000;
                 char22_0[  7] <= 32'h00000000;
                 char22_0[  8] <= 32'h00000000;
                 char22_0[  9] <= 32'h00000000;
                 char22_0[10] <= 32'h003FF000;
                 char22_0[11] <= 32'h00FFFC00;
                 char22_0[12] <= 32'h01F07E00;
                 char22_0[13] <= 32'h03C03F00;
                 char22_0[14] <= 32'h07801F80;
                 char22_0[15] <= 32'h0F800FC0;
                 char22_0[16] <= 32'h0F800FC0;
                 char22_0[17] <= 32'h0F8007E0;
                 char22_0[18] <= 32'h0FC007E0;
                 char22_0[19] <= 32'h0FC007E0;
                 char22_0[20] <= 32'h0FC007E0;
                 char22_0[21] <= 32'h07C007E0;
                 char22_0[22] <= 32'h000007E0;
                 char22_0[23] <= 32'h000007E0;
                 char22_0[24] <= 32'h000007C0;
                 char22_0[25] <= 32'h00000FC0;
                 char22_0[26] <= 32'h00000F80;
                 char22_0[27] <= 32'h00001F00;
                 char22_0[28] <= 32'h00007E00;
                 char22_0[29] <= 32'h0003FC00;
                 char22_0[30] <= 32'h001FF000;
                 char22_0[31] <= 32'h001FFC00;
                 char22_0[32] <= 32'h0000FF00;
                 char22_0[33] <= 32'h00001F80;
                 char22_0[34] <= 32'h00000FC0;
                 char22_0[35] <= 32'h000007E0;
                 char22_0[36] <= 32'h000003E0;
                 char22_0[37] <= 32'h000003F0;
                 char22_0[38] <= 32'h000003F0;
                 char22_0[39] <= 32'h000001F0;
                 char22_0[40] <= 32'h000001F8;
                 char22_0[41] <= 32'h000001F8;
                 char22_0[42] <= 32'h078001F8;
                 char22_0[43] <= 32'h0FC001F8;
                 char22_0[44] <= 32'h1FC001F8;
                 char22_0[45] <= 32'h1FC003F0;
                 char22_0[46] <= 32'h1FC003F0;
                 char22_0[47] <= 32'h1FC003E0;
                 char22_0[48] <= 32'h0F8007E0;
                 char22_0[49] <= 32'h0F8007C0;
                 char22_0[50] <= 32'h07C01F80;
                 char22_0[51] <= 32'h03F07F00;
                 char22_0[52] <= 32'h01FFFE00;
                 char22_0[53] <= 32'h003FF000;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//3
             4'd4: begin
                 char22_0[  0] <= 32'h00000000;
                 char22_0[  1] <= 32'h00000000;
                 char22_0[  2] <= 32'h00000000;
                 char22_0[  3] <= 32'h00000000;
                 char22_0[  4] <= 32'h00000000;
                 char22_0[  5] <= 32'h00000000;
                 char22_0[  6] <= 32'h00000000;
                 char22_0[  7] <= 32'h00000000;
                 char22_0[  8] <= 32'h00000000;
                 char22_0[  9] <= 32'h00000000;
                 char22_0[10] <= 32'h00001F00;
                 char22_0[11] <= 32'h00001F00;
                 char22_0[12] <= 32'h00003F00;
                 char22_0[13] <= 32'h00003F00;
                 char22_0[14] <= 32'h00007F00;
                 char22_0[15] <= 32'h0000FF00;
                 char22_0[16] <= 32'h0000FF00;
                 char22_0[17] <= 32'h0001FF00;
                 char22_0[18] <= 32'h0003FF00;
                 char22_0[19] <= 32'h0003BF00;
                 char22_0[20] <= 32'h0007BF00;
                 char22_0[21] <= 32'h00073F00;
                 char22_0[22] <= 32'h000F3F00;
                 char22_0[23] <= 32'h001E3F00;
                 char22_0[24] <= 32'h001C3F00;
                 char22_0[25] <= 32'h003C3F00;
                 char22_0[26] <= 32'h00783F00;
                 char22_0[27] <= 32'h00783F00;
                 char22_0[28] <= 32'h00F03F00;
                 char22_0[29] <= 32'h00E03F00;
                 char22_0[30] <= 32'h01E03F00;
                 char22_0[31] <= 32'h03C03F00;
                 char22_0[32] <= 32'h03803F00;
                 char22_0[33] <= 32'h07803F00;
                 char22_0[34] <= 32'h0F003F00;
                 char22_0[35] <= 32'h0F003F00;
                 char22_0[36] <= 32'h1E003F00;
                 char22_0[37] <= 32'h1C003F00;
                 char22_0[38] <= 32'h3C003F00;
                 char22_0[39] <= 32'h7FFFFFFE;
                 char22_0[40] <= 32'h7FFFFFFE;
                 char22_0[41] <= 32'h00003F00;
                 char22_0[42] <= 32'h00003F00;
                 char22_0[43] <= 32'h00003F00;
                 char22_0[44] <= 32'h00003F00;
                 char22_0[45] <= 32'h00003F00;
                 char22_0[46] <= 32'h00003F00;
                 char22_0[47] <= 32'h00003F00;
                 char22_0[48] <= 32'h00003F00;
                 char22_0[49] <= 32'h00003F00;
                 char22_0[50] <= 32'h00003F00;
                 char22_0[51] <= 32'h00007F80;
                 char22_0[52] <= 32'h000FFFFC;
                 char22_0[53] <= 32'h000FFFFC;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//4
             4'd5: begin
                 char22_0[  0] <= 32'h00000000;
                 char22_0[  1] <= 32'h00000000;
                 char22_0[  2] <= 32'h00000000;
                 char22_0[  3] <= 32'h00000000;
                 char22_0[  4] <= 32'h00000000;
                 char22_0[  5] <= 32'h00000000;
                 char22_0[  6] <= 32'h00000000;
                 char22_0[  7] <= 32'h00000000;
                 char22_0[  8] <= 32'h00000000;
                 char22_0[  9] <= 32'h00000000;
                 char22_0[10] <= 32'h00000000;
                 char22_0[11] <= 32'h03FFFFF0;
                 char22_0[12] <= 32'h03FFFFF0;
                 char22_0[13] <= 32'h03FFFFF0;
                 char22_0[14] <= 32'h03FFFFE0;
                 char22_0[15] <= 32'h03800000;
                 char22_0[16] <= 32'h03800000;
                 char22_0[17] <= 32'h03800000;
                 char22_0[18] <= 32'h03800000;
                 char22_0[19] <= 32'h03800000;
                 char22_0[20] <= 32'h07800000;
                 char22_0[21] <= 32'h07800000;
                 char22_0[22] <= 32'h07800000;
                 char22_0[23] <= 32'h07800000;
                 char22_0[24] <= 32'h07800000;
                 char22_0[25] <= 32'h07800000;
                 char22_0[26] <= 32'h078FF800;
                 char22_0[27] <= 32'h073FFE00;
                 char22_0[28] <= 32'h077FFF80;
                 char22_0[29] <= 32'h07FC3F80;
                 char22_0[30] <= 32'h07E00FC0;
                 char22_0[31] <= 32'h07C007E0;
                 char22_0[32] <= 32'h078007E0;
                 char22_0[33] <= 32'h078003F0;
                 char22_0[34] <= 32'h000003F0;
                 char22_0[35] <= 32'h000001F0;
                 char22_0[36] <= 32'h000001F8;
                 char22_0[37] <= 32'h000001F8;
                 char22_0[38] <= 32'h000001F8;
                 char22_0[39] <= 32'h000001F8;
                 char22_0[40] <= 32'h000001F8;
                 char22_0[41] <= 32'h078001F8;
                 char22_0[42] <= 32'h0FC001F8;
                 char22_0[43] <= 32'h1FC001F0;
                 char22_0[44] <= 32'h1FC001F0;
                 char22_0[45] <= 32'h1FC003F0;
                 char22_0[46] <= 32'h1F8003F0;
                 char22_0[47] <= 32'h1F8003E0;
                 char22_0[48] <= 32'h0F8007E0;
                 char22_0[49] <= 32'h078007C0;
                 char22_0[50] <= 32'h07C01F80;
                 char22_0[51] <= 32'h03F83F00;
                 char22_0[52] <= 32'h00FFFE00;
                 char22_0[53] <= 32'h003FF800;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//5
             4'd6: begin
                 char22_0[0] <= 32'h00000000;
                 char22_0[1] <= 32'h00000000;
                 char22_0[2] <= 32'h00000000;
                 char22_0[3] <= 32'h00000000;
                 char22_0[4] <= 32'h00000000;
                 char22_0[5] <= 32'h00000000;
                 char22_0[6] <= 32'h00000000;
                 char22_0[7] <= 32'h00000000;
                 char22_0[8] <= 32'h00000000;
                 char22_0[9] <= 32'h00000000;
                 char22_0[10] <= 32'h0007FE00;
                 char22_0[11] <= 32'h001FFF80;
                 char22_0[12] <= 32'h003F0FC0;
                 char22_0[13] <= 32'h007C07C0;
                 char22_0[14] <= 32'h00F807E0;
                 char22_0[15] <= 32'h01F007E0;
                 char22_0[16] <= 32'h03E007E0;
                 char22_0[17] <= 32'h03C007E0;
                 char22_0[18] <= 32'h07C003C0;
                 char22_0[19] <= 32'h07C00000;
                 char22_0[20] <= 32'h0FC00000;
                 char22_0[21] <= 32'h0F800000;
                 char22_0[22] <= 32'h0F800000;
                 char22_0[23] <= 32'h1F800000;
                 char22_0[24] <= 32'h1F800000;
                 char22_0[25] <= 32'h1F800000;
                 char22_0[26] <= 32'h1F87FE00;
                 char22_0[27] <= 32'h1F9FFF80;
                 char22_0[28] <= 32'h1FBFFFC0;
                 char22_0[29] <= 32'h3FFE1FC0;
                 char22_0[30] <= 32'h3FF807E0;
                 char22_0[31] <= 32'h3FE003F0;
                 char22_0[32] <= 32'h3FE003F0;
                 char22_0[33] <= 32'h3FC001F8;
                 char22_0[34] <= 32'h3F8001F8;
                 char22_0[35] <= 32'h3F8001F8;
                 char22_0[36] <= 32'h3F8000F8;
                 char22_0[37] <= 32'h3F8000F8;
                 char22_0[38] <= 32'h3F8000F8;
                 char22_0[39] <= 32'h1F8000F8;
                 char22_0[40] <= 32'h1F8000F8;
                 char22_0[41] <= 32'h1F8000F8;
                 char22_0[42] <= 32'h1F8000F8;
                 char22_0[43] <= 32'h1F8000F8;
                 char22_0[44] <= 32'h0FC001F8;
                 char22_0[45] <= 32'h0FC001F8;
                 char22_0[46] <= 32'h0FC001F0;
                 char22_0[47] <= 32'h07E001F0;
                 char22_0[48] <= 32'h03E003E0;
                 char22_0[49] <= 32'h03F003E0;
                 char22_0[50] <= 32'h01F807C0;
                 char22_0[51] <= 32'h00FE1F80;
                 char22_0[52] <= 32'h007FFE00;
                 char22_0[53] <= 32'h001FF800;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//6
             4'd7: begin
                 char22_0[0] <= 32'h00000000;
                 char22_0[1] <= 32'h00000000;
                 char22_0[2] <= 32'h00000000;
                 char22_0[3] <= 32'h00000000;
                 char22_0[4] <= 32'h00000000;
                 char22_0[5] <= 32'h00000000;
                 char22_0[6] <= 32'h00000000;
                 char22_0[7] <= 32'h00000000;
                 char22_0[8] <= 32'h00000000;
                 char22_0[9] <= 32'h00000000;
                 char22_0[10] <= 32'h00000000;
                 char22_0[11] <= 32'h07FFFFF8;
                 char22_0[12] <= 32'h07FFFFF8;
                 char22_0[13] <= 32'h07FFFFF8;
                 char22_0[14] <= 32'h0FFFFFF0;
                 char22_0[15] <= 32'h0FC000E0;
                 char22_0[16] <= 32'h0F8001E0;
                 char22_0[17] <= 32'h0F0001C0;
                 char22_0[18] <= 32'h0E0003C0;
                 char22_0[19] <= 32'h0E000780;
                 char22_0[20] <= 32'h1E000780;
                 char22_0[21] <= 32'h1C000F00;
                 char22_0[22] <= 32'h00000F00;
                 char22_0[23] <= 32'h00001E00;
                 char22_0[24] <= 32'h00001E00;
                 char22_0[25] <= 32'h00003C00;
                 char22_0[26] <= 32'h00003C00;
                 char22_0[27] <= 32'h00007800;
                 char22_0[28] <= 32'h00007800;
                 char22_0[29] <= 32'h0000F800;
                 char22_0[30] <= 32'h0000F000;
                 char22_0[31] <= 32'h0001F000;
                 char22_0[32] <= 32'h0001E000;
                 char22_0[33] <= 32'h0003E000;
                 char22_0[34] <= 32'h0003E000;
                 char22_0[35] <= 32'h0003E000;
                 char22_0[36] <= 32'h0007C000;
                 char22_0[37] <= 32'h0007C000;
                 char22_0[38] <= 32'h0007C000;
                 char22_0[39] <= 32'h000FC000;
                 char22_0[40] <= 32'h000FC000;
                 char22_0[41] <= 32'h000FC000;
                 char22_0[42] <= 32'h000FC000;
                 char22_0[43] <= 32'h001FC000;
                 char22_0[44] <= 32'h001FC000;
                 char22_0[45] <= 32'h001FC000;
                 char22_0[46] <= 32'h001FC000;
                 char22_0[47] <= 32'h001FC000;
                 char22_0[48] <= 32'h001FC000;
                 char22_0[49] <= 32'h001FC000;
                 char22_0[50] <= 32'h001FC000;
                 char22_0[51] <= 32'h001FC000;
                 char22_0[52] <= 32'h001FC000;
                 char22_0[53] <= 32'h000F8000;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//7
             4'd8: begin
                 char22_0[0] <= 32'h00000000;
                 char22_0[1] <= 32'h00000000;
                 char22_0[2] <= 32'h00000000;
                 char22_0[3] <= 32'h00000000;
                 char22_0[4] <= 32'h00000000;
                 char22_0[5] <= 32'h00000000;
                 char22_0[6] <= 32'h00000000;
                 char22_0[7] <= 32'h00000000;
                 char22_0[8] <= 32'h00000000;
                 char22_0[9] <= 32'h00000000;
                 char22_0[10] <= 32'h003FF800;
                 char22_0[11] <= 32'h00FFFE00;
                 char22_0[12] <= 32'h01F81F80;
                 char22_0[13] <= 32'h03E00FC0;
                 char22_0[14] <= 32'h07C003E0;
                 char22_0[15] <= 32'h0F8003E0;
                 char22_0[16] <= 32'h0F8001F0;
                 char22_0[17] <= 32'h1F0001F0;
                 char22_0[18] <= 32'h1F0001F0;
                 char22_0[19] <= 32'h1F0001F0;
                 char22_0[20] <= 32'h1F0001F0;
                 char22_0[21] <= 32'h1F0001F0;
                 char22_0[22] <= 32'h1F8001F0;
                 char22_0[23] <= 32'h1FC001F0;
                 char22_0[24] <= 32'h0FC001F0;
                 char22_0[25] <= 32'h0FF003E0;
                 char22_0[26] <= 32'h07F803C0;
                 char22_0[27] <= 32'h03FE0F80;
                 char22_0[28] <= 32'h01FF9F00;
                 char22_0[29] <= 32'h00FFFE00;
                 char22_0[30] <= 32'h003FF800;
                 char22_0[31] <= 32'h007FFC00;
                 char22_0[32] <= 32'h01F7FF00;
                 char22_0[33] <= 32'h03E1FF80;
                 char22_0[34] <= 32'h07C07FC0;
                 char22_0[35] <= 32'h0F801FE0;
                 char22_0[36] <= 32'h0F800FE0;
                 char22_0[37] <= 32'h1F0007F0;
                 char22_0[38] <= 32'h1F0003F0;
                 char22_0[39] <= 32'h3E0001F8;
                 char22_0[40] <= 32'h3E0001F8;
                 char22_0[41] <= 32'h3E0001F8;
                 char22_0[42] <= 32'h3E0000F8;
                 char22_0[43] <= 32'h3E0000F8;
                 char22_0[44] <= 32'h3E0000F8;
                 char22_0[45] <= 32'h3E0000F8;
                 char22_0[46] <= 32'h1F0001F0;
                 char22_0[47] <= 32'h1F0001F0;
                 char22_0[48] <= 32'h0F8003E0;
                 char22_0[49] <= 32'h0FC003E0;
                 char22_0[50] <= 32'h07E007C0;
                 char22_0[51] <= 32'h01F83F80;
                 char22_0[52] <= 32'h00FFFE00;
                 char22_0[53] <= 32'h003FF800;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//8
             4'd9: begin
                 char22_0[0] <= 32'h00000000;
                 char22_0[1] <= 32'h00000000;
                 char22_0[2] <= 32'h00000000;
                 char22_0[3] <= 32'h00000000;
                 char22_0[4] <= 32'h00000000;
                 char22_0[5] <= 32'h00000000;
                 char22_0[6] <= 32'h00000000;
                 char22_0[7] <= 32'h00000000;
                 char22_0[8] <= 32'h00000000;
                 char22_0[9] <= 32'h00000000;
                 char22_0[10] <= 32'h003FF000;
                 char22_0[11] <= 32'h00FFFC00;
                 char22_0[12] <= 32'h01F83F00;
                 char22_0[13] <= 32'h03E01F80;
                 char22_0[14] <= 32'h07C00F80;
                 char22_0[15] <= 32'h0FC007C0;
                 char22_0[16] <= 32'h0F8003E0;
                 char22_0[17] <= 32'h1F8003E0;
                 char22_0[18] <= 32'h1F0003F0;
                 char22_0[19] <= 32'h1F0003F0;
                 char22_0[20] <= 32'h3F0001F0;
                 char22_0[21] <= 32'h3F0001F0;
                 char22_0[22] <= 32'h3F0001F8;
                 char22_0[23] <= 32'h3F0001F8;
                 char22_0[24] <= 32'h3F0001F8;
                 char22_0[25] <= 32'h3F0001F8;
                 char22_0[26] <= 32'h3F0001F8;
                 char22_0[27] <= 32'h3F0001F8;
                 char22_0[28] <= 32'h3F0003F8;
                 char22_0[29] <= 32'h1F8003F8;
                 char22_0[30] <= 32'h1F8007F8;
                 char22_0[31] <= 32'h1F800FF8;
                 char22_0[32] <= 32'h0FC01FF8;
                 char22_0[33] <= 32'h0FE03FF8;
                 char22_0[34] <= 32'h07F8FDF8;
                 char22_0[35] <= 32'h03FFF9F8;
                 char22_0[36] <= 32'h01FFF1F8;
                 char22_0[37] <= 32'h003F83F8;
                 char22_0[38] <= 32'h000003F0;
                 char22_0[39] <= 32'h000003F0;
                 char22_0[40] <= 32'h000003F0;
                 char22_0[41] <= 32'h000003F0;
                 char22_0[42] <= 32'h000007E0;
                 char22_0[43] <= 32'h000007E0;
                 char22_0[44] <= 32'h000007C0;
                 char22_0[45] <= 32'h03C007C0;
                 char22_0[46] <= 32'h07C00F80;
                 char22_0[47] <= 32'h0FE00F80;
                 char22_0[48] <= 32'h0FE01F00;
                 char22_0[49] <= 32'h0FE03E00;
                 char22_0[50] <= 32'h07E07E00;
                 char22_0[51] <= 32'h07F1F800;
                 char22_0[52] <= 32'h03FFF000;
                 char22_0[53] <= 32'h00FFC000;
                 char22_0[54] <= 32'h00000000;
                 char22_0[55] <= 32'h00000000;
                 char22_0[56] <= 32'h00000000;
                 char22_0[57] <= 32'h00000000;
                 char22_0[58] <= 32'h00000000;
                 char22_0[59] <= 32'h00000000;
                 char22_0[60] <= 32'h00000000;
                 char22_0[61] <= 32'h00000000;
                 char22_0[62] <= 32'h00000000;
                 char22_0[63] <= 32'h00000000;
             end//9
             default: begin
                 char22_0[0] <= char22_0[0];
                 char22_0[1] <= char22_0[1];
                 char22_0[2] <= char22_0[2];
                 char22_0[3] <= char22_0[3];
                 char22_0[4] <= char22_0[4];
                 char22_0[5] <= char22_0[5];
                 char22_0[6] <= char22_0[6];
                 char22_0[7] <= char22_0[7];
                 char22_0[8] <= char22_0[8];
                 char22_0[9] <= char22_0[9];
                 char22_0[10] <= char22_0[10];
                 char22_0[11] <= char22_0[11];
                 char22_0[12] <= char22_0[12];
                 char22_0[13] <= char22_0[13];
                 char22_0[14] <= char22_0[14];
                 char22_0[15] <= char22_0[15];
                 char22_0[16] <= char22_0[16];
                 char22_0[17] <= char22_0[17];
                 char22_0[18] <= char22_0[18];
                 char22_0[19] <= char22_0[19];
                 char22_0[20] <= char22_0[20];
                 char22_0[21] <= char22_0[21];
                 char22_0[22] <= char22_0[22];
                 char22_0[23] <= char22_0[23];
                 char22_0[24] <= char22_0[24];
                 char22_0[25] <= char22_0[25];
                 char22_0[26] <= char22_0[26];
                 char22_0[27] <= char22_0[27];
                 char22_0[28] <= char22_0[28];
                 char22_0[29] <= char22_0[29];
                 char22_0[30] <= char22_0[30];
                 char22_0[31] <= char22_0[31];
                 char22_0[32] <= char22_0[32];
                 char22_0[33] <= char22_0[33];
                 char22_0[34] <= char22_0[34];
                 char22_0[35] <= char22_0[35];
                 char22_0[36] <= char22_0[36];
                 char22_0[37] <= char22_0[37];
                 char22_0[38] <= char22_0[38];
                 char22_0[39] <= char22_0[39];
                 char22_0[40] <= char22_0[40];
                 char22_0[41] <= char22_0[41];
                 char22_0[42] <= char22_0[42];
                 char22_0[43] <= char22_0[43];
                 char22_0[44] <= char22_0[44];
                 char22_0[45] <= char22_0[45];
                 char22_0[46] <= char22_0[46];
                 char22_0[47] <= char22_0[47];
                 char22_0[48] <= char22_0[48];
                 char22_0[49] <= char22_0[49];
                 char22_0[50] <= char22_0[50];
                 char22_0[51] <= char22_0[51];
                 char22_0[52] <= char22_0[52];
                 char22_0[53] <= char22_0[53];
                 char22_0[54] <= char22_0[54];
                 char22_0[55] <= char22_0[55];
                 char22_0[56] <= char22_0[56];
                 char22_0[57] <= char22_0[57];
                 char22_0[58] <= char22_0[58];
                 char22_0[59] <= char22_0[59];
                 char22_0[60] <= char22_0[60];
                 char22_0[61] <= char22_0[61];
                 char22_0[62] <= char22_0[62];
                 char22_0[63] <= char22_0[63];
             end
         endcase
     
         case((li - hkm*(li/hkm))/tenkm)
                 4'd0: begin
                     char22_1[  0] <= 32'h00000000;
                     char22_1[  1] <= 32'h00000000;
                     char22_1[  2] <= 32'h00000000;
                     char22_1[  3] <= 32'h00000000;
                     char22_1[  4] <= 32'h00000000;
                     char22_1[  5] <= 32'h00000000;
                     char22_1[  6] <= 32'h00000000;
                     char22_1[  7] <= 32'h00000000;
                     char22_1[  8] <= 32'h00000000;
                     char22_1[  9] <= 32'h00000000;
                     char22_1[10] <= 32'h000FF000;
                     char22_1[11] <= 32'h003FFC00;
                     char22_1[12] <= 32'h007E7E00;
                     char22_1[13] <= 32'h00F81F00;
                     char22_1[14] <= 32'h01F00F80;
                     char22_1[15] <= 32'h03F00FC0;
                     char22_1[16] <= 32'h03E007C0;
                     char22_1[17] <= 32'h07E007E0;
                     char22_1[18] <= 32'h07C003E0;
                     char22_1[19] <= 32'h0FC003F0;
                     char22_1[20] <= 32'h0FC003F0;
                     char22_1[21] <= 32'h0FC003F0;
                     char22_1[22] <= 32'h1F8001F8;
                     char22_1[23] <= 32'h1F8001F8;
                     char22_1[24] <= 32'h1F8001F8;
                     char22_1[25] <= 32'h1F8001F8;
                     char22_1[26] <= 32'h1F8001F8;
                     char22_1[27] <= 32'h3F8001F8;
                     char22_1[28] <= 32'h3F8001F8;
                     char22_1[29] <= 32'h3F8001F8;
                     char22_1[30] <= 32'h3F8001F8;
                     char22_1[31] <= 32'h3F8001F8;
                     char22_1[32] <= 32'h3F8001F8;
                     char22_1[33] <= 32'h3F8001F8;
                     char22_1[34] <= 32'h3F8001F8;
                     char22_1[35] <= 32'h3F8001F8;
                     char22_1[36] <= 32'h3F8001F8;
                     char22_1[37] <= 32'h1F8001F8;
                     char22_1[38] <= 32'h1F8001F8;
                     char22_1[39] <= 32'h1F8001F8;
                     char22_1[40] <= 32'h1F8001F8;
                     char22_1[41] <= 32'h1F8001F0;
                     char22_1[42] <= 32'h0F8003F0;
                     char22_1[43] <= 32'h0FC003F0;
                     char22_1[44] <= 32'h0FC003F0;
                     char22_1[45] <= 32'h07C003E0;
                     char22_1[46] <= 32'h07E007E0;
                     char22_1[47] <= 32'h03E007C0;
                     char22_1[48] <= 32'h03F00FC0;
                     char22_1[49] <= 32'h01F00F80;
                     char22_1[50] <= 32'h00F81F00;
                     char22_1[51] <= 32'h007E7E00;
                     char22_1[52] <= 32'h003FFC00;
                     char22_1[53] <= 32'h000FF000;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//0
                 4'd1: begin
                     char22_1[  0] <= 32'h00000000;
                     char22_1[  1] <= 32'h00000000;
                     char22_1[  2] <= 32'h00000000;
                     char22_1[  3] <= 32'h00000000;
                     char22_1[  4] <= 32'h00000000;
                     char22_1[  5] <= 32'h00000000;
                     char22_1[  6] <= 32'h00000000;
                     char22_1[  7] <= 32'h00000000;
                     char22_1[  8] <= 32'h00000000;
                     char22_1[  9] <= 32'h00000000;
                     char22_1[10] <= 32'h0000E000;
                     char22_1[11] <= 32'h0001E000;
                     char22_1[12] <= 32'h0003E000;
                     char22_1[13] <= 32'h001FE000;
                     char22_1[14] <= 32'h03FFE000;
                     char22_1[15] <= 32'h03FFE000;
                     char22_1[16] <= 32'h0007E000;
                     char22_1[17] <= 32'h0007E000;
                     char22_1[18] <= 32'h0007E000;
                     char22_1[19] <= 32'h0007E000;
                     char22_1[20] <= 32'h0007E000;
                     char22_1[21] <= 32'h0007E000;
                     char22_1[22] <= 32'h0007E000;
                     char22_1[23] <= 32'h0007E000;
                     char22_1[24] <= 32'h0007E000;
                     char22_1[25] <= 32'h0007E000;
                     char22_1[26] <= 32'h0007E000;
                     char22_1[27] <= 32'h0007E000;
                     char22_1[28] <= 32'h0007E000;
                     char22_1[29] <= 32'h0007E000;
                     char22_1[30] <= 32'h0007E000;
                     char22_1[31] <= 32'h0007E000;
                     char22_1[32] <= 32'h0007E000;
                     char22_1[33] <= 32'h0007E000;
                     char22_1[34] <= 32'h0007E000;
                     char22_1[35] <= 32'h0007E000;
                     char22_1[36] <= 32'h0007E000;
                     char22_1[37] <= 32'h0007E000;
                     char22_1[38] <= 32'h0007E000;
                     char22_1[39] <= 32'h0007E000;
                     char22_1[40] <= 32'h0007E000;
                     char22_1[41] <= 32'h0007E000;
                     char22_1[42] <= 32'h0007E000;
                     char22_1[43] <= 32'h0007E000;
                     char22_1[44] <= 32'h0007E000;
                     char22_1[45] <= 32'h0007E000;
                     char22_1[46] <= 32'h0007E000;
                     char22_1[47] <= 32'h0007E000;
                     char22_1[48] <= 32'h0007E000;
                     char22_1[49] <= 32'h0007E000;
                     char22_1[50] <= 32'h0007E000;
                     char22_1[51] <= 32'h000FF800;
                     char22_1[52] <= 32'h03FFFFC0;
                     char22_1[53] <= 32'h03FFFFC0;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//1
                 4'd2: begin
                     char22_1[  0] <= 32'h00000000;
                     char22_1[  1] <= 32'h00000000;
                     char22_1[  2] <= 32'h00000000;
                     char22_1[  3] <= 32'h00000000;
                     char22_1[  4] <= 32'h00000000;
                     char22_1[  5] <= 32'h00000000;
                     char22_1[  6] <= 32'h00000000;
                     char22_1[  7] <= 32'h00000000;
                     char22_1[  8] <= 32'h00000000;
                     char22_1[  9] <= 32'h00000000;
                     char22_1[10] <= 32'h001FFC00;
                     char22_1[11] <= 32'h007FFF00;
                     char22_1[12] <= 32'h01F83F80;
                     char22_1[13] <= 32'h03E00FC0;
                     char22_1[14] <= 32'h07C007E0;
                     char22_1[15] <= 32'h078007E0;
                     char22_1[16] <= 32'h0F8003F0;
                     char22_1[17] <= 32'h0F8003F0;
                     char22_1[18] <= 32'h1F8003F0;
                     char22_1[19] <= 32'h1F8003F0;
                     char22_1[20] <= 32'h1FC003F0;
                     char22_1[21] <= 32'h1FC003F0;
                     char22_1[22] <= 32'h1FC003F0;
                     char22_1[23] <= 32'h0FC003F0;
                     char22_1[24] <= 32'h07C003F0;
                     char22_1[25] <= 32'h000003E0;
                     char22_1[26] <= 32'h000007E0;
                     char22_1[27] <= 32'h000007E0;
                     char22_1[28] <= 32'h00000FC0;
                     char22_1[29] <= 32'h00000F80;
                     char22_1[30] <= 32'h00001F80;
                     char22_1[31] <= 32'h00003F00;
                     char22_1[32] <= 32'h00003E00;
                     char22_1[33] <= 32'h00007C00;
                     char22_1[34] <= 32'h0000F800;
                     char22_1[35] <= 32'h0001F000;
                     char22_1[36] <= 32'h0003E000;
                     char22_1[37] <= 32'h0007C000;
                     char22_1[38] <= 32'h000F8000;
                     char22_1[39] <= 32'h001F0000;
                     char22_1[40] <= 32'h003E0000;
                     char22_1[41] <= 32'h007C0000;
                     char22_1[42] <= 32'h00F80000;
                     char22_1[43] <= 32'h01F00038;
                     char22_1[44] <= 32'h01E00038;
                     char22_1[45] <= 32'h03C00070;
                     char22_1[46] <= 32'h07800070;
                     char22_1[47] <= 32'h0F8000F0;
                     char22_1[48] <= 32'h0F0000F0;
                     char22_1[49] <= 32'h1E0003F0;
                     char22_1[50] <= 32'h3FFFFFF0;
                     char22_1[51] <= 32'h3FFFFFF0;
                     char22_1[52] <= 32'h3FFFFFE0;
                     char22_1[53] <= 32'h3FFFFFE0;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//2
                 4'd3: begin
                     char22_1[  0] <= 32'h00000000;
                     char22_1[  1] <= 32'h00000000;
                     char22_1[  2] <= 32'h00000000;
                     char22_1[  3] <= 32'h00000000;
                     char22_1[  4] <= 32'h00000000;
                     char22_1[  5] <= 32'h00000000;
                     char22_1[  6] <= 32'h00000000;
                     char22_1[  7] <= 32'h00000000;
                     char22_1[  8] <= 32'h00000000;
                     char22_1[  9] <= 32'h00000000;
                     char22_1[10] <= 32'h003FF000;
                     char22_1[11] <= 32'h00FFFC00;
                     char22_1[12] <= 32'h01F07E00;
                     char22_1[13] <= 32'h03C03F00;
                     char22_1[14] <= 32'h07801F80;
                     char22_1[15] <= 32'h0F800FC0;
                     char22_1[16] <= 32'h0F800FC0;
                     char22_1[17] <= 32'h0F8007E0;
                     char22_1[18] <= 32'h0FC007E0;
                     char22_1[19] <= 32'h0FC007E0;
                     char22_1[20] <= 32'h0FC007E0;
                     char22_1[21] <= 32'h07C007E0;
                     char22_1[22] <= 32'h000007E0;
                     char22_1[23] <= 32'h000007E0;
                     char22_1[24] <= 32'h000007C0;
                     char22_1[25] <= 32'h00000FC0;
                     char22_1[26] <= 32'h00000F80;
                     char22_1[27] <= 32'h00001F00;
                     char22_1[28] <= 32'h00007E00;
                     char22_1[29] <= 32'h0003FC00;
                     char22_1[30] <= 32'h001FF000;
                     char22_1[31] <= 32'h001FFC00;
                     char22_1[32] <= 32'h0000FF00;
                     char22_1[33] <= 32'h00001F80;
                     char22_1[34] <= 32'h00000FC0;
                     char22_1[35] <= 32'h000007E0;
                     char22_1[36] <= 32'h000003E0;
                     char22_1[37] <= 32'h000003F0;
                     char22_1[38] <= 32'h000003F0;
                     char22_1[39] <= 32'h000001F0;
                     char22_1[40] <= 32'h000001F8;
                     char22_1[41] <= 32'h000001F8;
                     char22_1[42] <= 32'h078001F8;
                     char22_1[43] <= 32'h0FC001F8;
                     char22_1[44] <= 32'h1FC001F8;
                     char22_1[45] <= 32'h1FC003F0;
                     char22_1[46] <= 32'h1FC003F0;
                     char22_1[47] <= 32'h1FC003E0;
                     char22_1[48] <= 32'h0F8007E0;
                     char22_1[49] <= 32'h0F8007C0;
                     char22_1[50] <= 32'h07C01F80;
                     char22_1[51] <= 32'h03F07F00;
                     char22_1[52] <= 32'h01FFFE00;
                     char22_1[53] <= 32'h003FF000;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//3
                 4'd4: begin
                     char22_1[  0] <= 32'h00000000;
                     char22_1[  1] <= 32'h00000000;
                     char22_1[  2] <= 32'h00000000;
                     char22_1[  3] <= 32'h00000000;
                     char22_1[  4] <= 32'h00000000;
                     char22_1[  5] <= 32'h00000000;
                     char22_1[  6] <= 32'h00000000;
                     char22_1[  7] <= 32'h00000000;
                     char22_1[  8] <= 32'h00000000;
                     char22_1[  9] <= 32'h00000000;
                     char22_1[10] <= 32'h00001F00;
                     char22_1[11] <= 32'h00001F00;
                     char22_1[12] <= 32'h00003F00;
                     char22_1[13] <= 32'h00003F00;
                     char22_1[14] <= 32'h00007F00;
                     char22_1[15] <= 32'h0000FF00;
                     char22_1[16] <= 32'h0000FF00;
                     char22_1[17] <= 32'h0001FF00;
                     char22_1[18] <= 32'h0003FF00;
                     char22_1[19] <= 32'h0003BF00;
                     char22_1[20] <= 32'h0007BF00;
                     char22_1[21] <= 32'h00073F00;
                     char22_1[22] <= 32'h000F3F00;
                     char22_1[23] <= 32'h001E3F00;
                     char22_1[24] <= 32'h001C3F00;
                     char22_1[25] <= 32'h003C3F00;
                     char22_1[26] <= 32'h00783F00;
                     char22_1[27] <= 32'h00783F00;
                     char22_1[28] <= 32'h00F03F00;
                     char22_1[29] <= 32'h00E03F00;
                     char22_1[30] <= 32'h01E03F00;
                     char22_1[31] <= 32'h03C03F00;
                     char22_1[32] <= 32'h03803F00;
                     char22_1[33] <= 32'h07803F00;
                     char22_1[34] <= 32'h0F003F00;
                     char22_1[35] <= 32'h0F003F00;
                     char22_1[36] <= 32'h1E003F00;
                     char22_1[37] <= 32'h1C003F00;
                     char22_1[38] <= 32'h3C003F00;
                     char22_1[39] <= 32'h7FFFFFFE;
                     char22_1[40] <= 32'h7FFFFFFE;
                     char22_1[41] <= 32'h00003F00;
                     char22_1[42] <= 32'h00003F00;
                     char22_1[43] <= 32'h00003F00;
                     char22_1[44] <= 32'h00003F00;
                     char22_1[45] <= 32'h00003F00;
                     char22_1[46] <= 32'h00003F00;
                     char22_1[47] <= 32'h00003F00;
                     char22_1[48] <= 32'h00003F00;
                     char22_1[49] <= 32'h00003F00;
                     char22_1[50] <= 32'h00003F00;
                     char22_1[51] <= 32'h00007F80;
                     char22_1[52] <= 32'h000FFFFC;
                     char22_1[53] <= 32'h000FFFFC;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//4
                 4'd5: begin
                     char22_1[  0] <= 32'h00000000;
                     char22_1[  1] <= 32'h00000000;
                     char22_1[  2] <= 32'h00000000;
                     char22_1[  3] <= 32'h00000000;
                     char22_1[  4] <= 32'h00000000;
                     char22_1[  5] <= 32'h00000000;
                     char22_1[  6] <= 32'h00000000;
                     char22_1[  7] <= 32'h00000000;
                     char22_1[  8] <= 32'h00000000;
                     char22_1[  9] <= 32'h00000000;
                     char22_1[10] <= 32'h00000000;
                     char22_1[11] <= 32'h03FFFFF0;
                     char22_1[12] <= 32'h03FFFFF0;
                     char22_1[13] <= 32'h03FFFFF0;
                     char22_1[14] <= 32'h03FFFFE0;
                     char22_1[15] <= 32'h03800000;
                     char22_1[16] <= 32'h03800000;
                     char22_1[17] <= 32'h03800000;
                     char22_1[18] <= 32'h03800000;
                     char22_1[19] <= 32'h03800000;
                     char22_1[20] <= 32'h07800000;
                     char22_1[21] <= 32'h07800000;
                     char22_1[22] <= 32'h07800000;
                     char22_1[23] <= 32'h07800000;
                     char22_1[24] <= 32'h07800000;
                     char22_1[25] <= 32'h07800000;
                     char22_1[26] <= 32'h078FF800;
                     char22_1[27] <= 32'h073FFE00;
                     char22_1[28] <= 32'h077FFF80;
                     char22_1[29] <= 32'h07FC3F80;
                     char22_1[30] <= 32'h07E00FC0;
                     char22_1[31] <= 32'h07C007E0;
                     char22_1[32] <= 32'h078007E0;
                     char22_1[33] <= 32'h078003F0;
                     char22_1[34] <= 32'h000003F0;
                     char22_1[35] <= 32'h000001F0;
                     char22_1[36] <= 32'h000001F8;
                     char22_1[37] <= 32'h000001F8;
                     char22_1[38] <= 32'h000001F8;
                     char22_1[39] <= 32'h000001F8;
                     char22_1[40] <= 32'h000001F8;
                     char22_1[41] <= 32'h078001F8;
                     char22_1[42] <= 32'h0FC001F8;
                     char22_1[43] <= 32'h1FC001F0;
                     char22_1[44] <= 32'h1FC001F0;
                     char22_1[45] <= 32'h1FC003F0;
                     char22_1[46] <= 32'h1F8003F0;
                     char22_1[47] <= 32'h1F8003E0;
                     char22_1[48] <= 32'h0F8007E0;
                     char22_1[49] <= 32'h078007C0;
                     char22_1[50] <= 32'h07C01F80;
                     char22_1[51] <= 32'h03F83F00;
                     char22_1[52] <= 32'h00FFFE00;
                     char22_1[53] <= 32'h003FF800;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//5
                 4'd6: begin
                     char22_1[0] <= 32'h00000000;
                     char22_1[1] <= 32'h00000000;
                     char22_1[2] <= 32'h00000000;
                     char22_1[3] <= 32'h00000000;
                     char22_1[4] <= 32'h00000000;
                     char22_1[5] <= 32'h00000000;
                     char22_1[6] <= 32'h00000000;
                     char22_1[7] <= 32'h00000000;
                     char22_1[8] <= 32'h00000000;
                     char22_1[9] <= 32'h00000000;
                     char22_1[10] <= 32'h0007FE00;
                     char22_1[11] <= 32'h001FFF80;
                     char22_1[12] <= 32'h003F0FC0;
                     char22_1[13] <= 32'h007C07C0;
                     char22_1[14] <= 32'h00F807E0;
                     char22_1[15] <= 32'h01F007E0;
                     char22_1[16] <= 32'h03E007E0;
                     char22_1[17] <= 32'h03C007E0;
                     char22_1[18] <= 32'h07C003C0;
                     char22_1[19] <= 32'h07C00000;
                     char22_1[20] <= 32'h0FC00000;
                     char22_1[21] <= 32'h0F800000;
                     char22_1[22] <= 32'h0F800000;
                     char22_1[23] <= 32'h1F800000;
                     char22_1[24] <= 32'h1F800000;
                     char22_1[25] <= 32'h1F800000;
                     char22_1[26] <= 32'h1F87FE00;
                     char22_1[27] <= 32'h1F9FFF80;
                     char22_1[28] <= 32'h1FBFFFC0;
                     char22_1[29] <= 32'h3FFE1FC0;
                     char22_1[30] <= 32'h3FF807E0;
                     char22_1[31] <= 32'h3FE003F0;
                     char22_1[32] <= 32'h3FE003F0;
                     char22_1[33] <= 32'h3FC001F8;
                     char22_1[34] <= 32'h3F8001F8;
                     char22_1[35] <= 32'h3F8001F8;
                     char22_1[36] <= 32'h3F8000F8;
                     char22_1[37] <= 32'h3F8000F8;
                     char22_1[38] <= 32'h3F8000F8;
                     char22_1[39] <= 32'h1F8000F8;
                     char22_1[40] <= 32'h1F8000F8;
                     char22_1[41] <= 32'h1F8000F8;
                     char22_1[42] <= 32'h1F8000F8;
                     char22_1[43] <= 32'h1F8000F8;
                     char22_1[44] <= 32'h0FC001F8;
                     char22_1[45] <= 32'h0FC001F8;
                     char22_1[46] <= 32'h0FC001F0;
                     char22_1[47] <= 32'h07E001F0;
                     char22_1[48] <= 32'h03E003E0;
                     char22_1[49] <= 32'h03F003E0;
                     char22_1[50] <= 32'h01F807C0;
                     char22_1[51] <= 32'h00FE1F80;
                     char22_1[52] <= 32'h007FFE00;
                     char22_1[53] <= 32'h001FF800;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//6
                 4'd7: begin
                     char22_1[0] <= 32'h00000000;
                     char22_1[1] <= 32'h00000000;
                     char22_1[2] <= 32'h00000000;
                     char22_1[3] <= 32'h00000000;
                     char22_1[4] <= 32'h00000000;
                     char22_1[5] <= 32'h00000000;
                     char22_1[6] <= 32'h00000000;
                     char22_1[7] <= 32'h00000000;
                     char22_1[8] <= 32'h00000000;
                     char22_1[9] <= 32'h00000000;
                     char22_1[10] <= 32'h00000000;
                     char22_1[11] <= 32'h07FFFFF8;
                     char22_1[12] <= 32'h07FFFFF8;
                     char22_1[13] <= 32'h07FFFFF8;
                     char22_1[14] <= 32'h0FFFFFF0;
                     char22_1[15] <= 32'h0FC000E0;
                     char22_1[16] <= 32'h0F8001E0;
                     char22_1[17] <= 32'h0F0001C0;
                     char22_1[18] <= 32'h0E0003C0;
                     char22_1[19] <= 32'h0E000780;
                     char22_1[20] <= 32'h1E000780;
                     char22_1[21] <= 32'h1C000F00;
                     char22_1[22] <= 32'h00000F00;
                     char22_1[23] <= 32'h00001E00;
                     char22_1[24] <= 32'h00001E00;
                     char22_1[25] <= 32'h00003C00;
                     char22_1[26] <= 32'h00003C00;
                     char22_1[27] <= 32'h00007800;
                     char22_1[28] <= 32'h00007800;
                     char22_1[29] <= 32'h0000F800;
                     char22_1[30] <= 32'h0000F000;
                     char22_1[31] <= 32'h0001F000;
                     char22_1[32] <= 32'h0001E000;
                     char22_1[33] <= 32'h0003E000;
                     char22_1[34] <= 32'h0003E000;
                     char22_1[35] <= 32'h0003E000;
                     char22_1[36] <= 32'h0007C000;
                     char22_1[37] <= 32'h0007C000;
                     char22_1[38] <= 32'h0007C000;
                     char22_1[39] <= 32'h000FC000;
                     char22_1[40] <= 32'h000FC000;
                     char22_1[41] <= 32'h000FC000;
                     char22_1[42] <= 32'h000FC000;
                     char22_1[43] <= 32'h001FC000;
                     char22_1[44] <= 32'h001FC000;
                     char22_1[45] <= 32'h001FC000;
                     char22_1[46] <= 32'h001FC000;
                     char22_1[47] <= 32'h001FC000;
                     char22_1[48] <= 32'h001FC000;
                     char22_1[49] <= 32'h001FC000;
                     char22_1[50] <= 32'h001FC000;
                     char22_1[51] <= 32'h001FC000;
                     char22_1[52] <= 32'h001FC000;
                     char22_1[53] <= 32'h000F8000;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//7
                 4'd8: begin
                     char22_1[0] <= 32'h00000000;
                     char22_1[1] <= 32'h00000000;
                     char22_1[2] <= 32'h00000000;
                     char22_1[3] <= 32'h00000000;
                     char22_1[4] <= 32'h00000000;
                     char22_1[5] <= 32'h00000000;
                     char22_1[6] <= 32'h00000000;
                     char22_1[7] <= 32'h00000000;
                     char22_1[8] <= 32'h00000000;
                     char22_1[9] <= 32'h00000000;
                     char22_1[10] <= 32'h003FF800;
                     char22_1[11] <= 32'h00FFFE00;
                     char22_1[12] <= 32'h01F81F80;
                     char22_1[13] <= 32'h03E00FC0;
                     char22_1[14] <= 32'h07C003E0;
                     char22_1[15] <= 32'h0F8003E0;
                     char22_1[16] <= 32'h0F8001F0;
                     char22_1[17] <= 32'h1F0001F0;
                     char22_1[18] <= 32'h1F0001F0;
                     char22_1[19] <= 32'h1F0001F0;
                     char22_1[20] <= 32'h1F0001F0;
                     char22_1[21] <= 32'h1F0001F0;
                     char22_1[22] <= 32'h1F8001F0;
                     char22_1[23] <= 32'h1FC001F0;
                     char22_1[24] <= 32'h0FC001F0;
                     char22_1[25] <= 32'h0FF003E0;
                     char22_1[26] <= 32'h07F803C0;
                     char22_1[27] <= 32'h03FE0F80;
                     char22_1[28] <= 32'h01FF9F00;
                     char22_1[29] <= 32'h00FFFE00;
                     char22_1[30] <= 32'h003FF800;
                     char22_1[31] <= 32'h007FFC00;
                     char22_1[32] <= 32'h01F7FF00;
                     char22_1[33] <= 32'h03E1FF80;
                     char22_1[34] <= 32'h07C07FC0;
                     char22_1[35] <= 32'h0F801FE0;
                     char22_1[36] <= 32'h0F800FE0;
                     char22_1[37] <= 32'h1F0007F0;
                     char22_1[38] <= 32'h1F0003F0;
                     char22_1[39] <= 32'h3E0001F8;
                     char22_1[40] <= 32'h3E0001F8;
                     char22_1[41] <= 32'h3E0001F8;
                     char22_1[42] <= 32'h3E0000F8;
                     char22_1[43] <= 32'h3E0000F8;
                     char22_1[44] <= 32'h3E0000F8;
                     char22_1[45] <= 32'h3E0000F8;
                     char22_1[46] <= 32'h1F0001F0;
                     char22_1[47] <= 32'h1F0001F0;
                     char22_1[48] <= 32'h0F8003E0;
                     char22_1[49] <= 32'h0FC003E0;
                     char22_1[50] <= 32'h07E007C0;
                     char22_1[51] <= 32'h01F83F80;
                     char22_1[52] <= 32'h00FFFE00;
                     char22_1[53] <= 32'h003FF800;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//8
                 4'd9: begin
                     char22_1[0] <= 32'h00000000;
                     char22_1[1] <= 32'h00000000;
                     char22_1[2] <= 32'h00000000;
                     char22_1[3] <= 32'h00000000;
                     char22_1[4] <= 32'h00000000;
                     char22_1[5] <= 32'h00000000;
                     char22_1[6] <= 32'h00000000;
                     char22_1[7] <= 32'h00000000;
                     char22_1[8] <= 32'h00000000;
                     char22_1[9] <= 32'h00000000;
                     char22_1[10] <= 32'h003FF000;
                     char22_1[11] <= 32'h00FFFC00;
                     char22_1[12] <= 32'h01F83F00;
                     char22_1[13] <= 32'h03E01F80;
                     char22_1[14] <= 32'h07C00F80;
                     char22_1[15] <= 32'h0FC007C0;
                     char22_1[16] <= 32'h0F8003E0;
                     char22_1[17] <= 32'h1F8003E0;
                     char22_1[18] <= 32'h1F0003F0;
                     char22_1[19] <= 32'h1F0003F0;
                     char22_1[20] <= 32'h3F0001F0;
                     char22_1[21] <= 32'h3F0001F0;
                     char22_1[22] <= 32'h3F0001F8;
                     char22_1[23] <= 32'h3F0001F8;
                     char22_1[24] <= 32'h3F0001F8;
                     char22_1[25] <= 32'h3F0001F8;
                     char22_1[26] <= 32'h3F0001F8;
                     char22_1[27] <= 32'h3F0001F8;
                     char22_1[28] <= 32'h3F0003F8;
                     char22_1[29] <= 32'h1F8003F8;
                     char22_1[30] <= 32'h1F8007F8;
                     char22_1[31] <= 32'h1F800FF8;
                     char22_1[32] <= 32'h0FC01FF8;
                     char22_1[33] <= 32'h0FE03FF8;
                     char22_1[34] <= 32'h07F8FDF8;
                     char22_1[35] <= 32'h03FFF9F8;
                     char22_1[36] <= 32'h01FFF1F8;
                     char22_1[37] <= 32'h003F83F8;
                     char22_1[38] <= 32'h000003F0;
                     char22_1[39] <= 32'h000003F0;
                     char22_1[40] <= 32'h000003F0;
                     char22_1[41] <= 32'h000003F0;
                     char22_1[42] <= 32'h000007E0;
                     char22_1[43] <= 32'h000007E0;
                     char22_1[44] <= 32'h000007C0;
                     char22_1[45] <= 32'h03C007C0;
                     char22_1[46] <= 32'h07C00F80;
                     char22_1[47] <= 32'h0FE00F80;
                     char22_1[48] <= 32'h0FE01F00;
                     char22_1[49] <= 32'h0FE03E00;
                     char22_1[50] <= 32'h07E07E00;
                     char22_1[51] <= 32'h07F1F800;
                     char22_1[52] <= 32'h03FFF000;
                     char22_1[53] <= 32'h00FFC000;
                     char22_1[54] <= 32'h00000000;
                     char22_1[55] <= 32'h00000000;
                     char22_1[56] <= 32'h00000000;
                     char22_1[57] <= 32'h00000000;
                     char22_1[58] <= 32'h00000000;
                     char22_1[59] <= 32'h00000000;
                     char22_1[60] <= 32'h00000000;
                     char22_1[61] <= 32'h00000000;
                     char22_1[62] <= 32'h00000000;
                     char22_1[63] <= 32'h00000000;
                 end//9
                 default: begin
                     char22_1[0] <= char22_1[0];
                     char22_1[1] <= char22_1[1];
                     char22_1[2] <= char22_1[2];
                     char22_1[3] <= char22_1[3];
                     char22_1[4] <= char22_1[4];
                     char22_1[5] <= char22_1[5];
                     char22_1[6] <= char22_1[6];
                     char22_1[7] <= char22_1[7];
                     char22_1[8] <= char22_1[8];
                     char22_1[9] <= char22_1[9];
                     char22_1[10] <= char22_1[10];
                     char22_1[11] <= char22_1[11];
                     char22_1[12] <= char22_1[12];
                     char22_1[13] <= char22_1[13];
                     char22_1[14] <= char22_1[14];
                     char22_1[15] <= char22_1[15];
                     char22_1[16] <= char22_1[16];
                     char22_1[17] <= char22_1[17];
                     char22_1[18] <= char22_1[18];
                     char22_1[19] <= char22_1[19];
                     char22_1[20] <= char22_1[20];
                     char22_1[21] <= char22_1[21];
                     char22_1[22] <= char22_1[22];
                     char22_1[23] <= char22_1[23];
                     char22_1[24] <= char22_1[24];
                     char22_1[25] <= char22_1[25];
                     char22_1[26] <= char22_1[26];
                     char22_1[27] <= char22_1[27];
                     char22_1[28] <= char22_1[28];
                     char22_1[29] <= char22_1[29];
                     char22_1[30] <= char22_1[30];
                     char22_1[31] <= char22_1[31];
                     char22_1[32] <= char22_1[32];
                     char22_1[33] <= char22_1[33];
                     char22_1[34] <= char22_1[34];
                     char22_1[35] <= char22_1[35];
                     char22_1[36] <= char22_1[36];
                     char22_1[37] <= char22_1[37];
                     char22_1[38] <= char22_1[38];
                     char22_1[39] <= char22_1[39];
                     char22_1[40] <= char22_1[40];
                     char22_1[41] <= char22_1[41];
                     char22_1[42] <= char22_1[42];
                     char22_1[43] <= char22_1[43];
                     char22_1[44] <= char22_1[44];
                     char22_1[45] <= char22_1[45];
                     char22_1[46] <= char22_1[46];
                     char22_1[47] <= char22_1[47];
                     char22_1[48] <= char22_1[48];
                     char22_1[49] <= char22_1[49];
                     char22_1[50] <= char22_1[50];
                     char22_1[51] <= char22_1[51];
                     char22_1[52] <= char22_1[52];
                     char22_1[53] <= char22_1[53];
                     char22_1[54] <= char22_1[54];
                     char22_1[55] <= char22_1[55];
                     char22_1[56] <= char22_1[56];
                     char22_1[57] <= char22_1[57];
                     char22_1[58] <= char22_1[58];
                     char22_1[59] <= char22_1[59];
                     char22_1[60] <= char22_1[60];
                     char22_1[61] <= char22_1[61];
                     char22_1[62] <= char22_1[62];
                     char22_1[63] <= char22_1[63];
                 end
             endcase
     
         case((li - tenkm*(li/tenkm))/onekm)
                 4'd0: begin
                     char22_2[  0] <= 32'h00000000;
                     char22_2[  1] <= 32'h00000000;
                     char22_2[  2] <= 32'h00000000;
                     char22_2[  3] <= 32'h00000000;
                     char22_2[  4] <= 32'h00000000;
                     char22_2[  5] <= 32'h00000000;
                     char22_2[  6] <= 32'h00000000;
                     char22_2[  7] <= 32'h00000000;
                     char22_2[  8] <= 32'h00000000;
                     char22_2[  9] <= 32'h00000000;
                     char22_2[10] <= 32'h000FF000;
                     char22_2[11] <= 32'h003FFC00;
                     char22_2[12] <= 32'h007E7E00;
                     char22_2[13] <= 32'h00F81F00;
                     char22_2[14] <= 32'h01F00F80;
                     char22_2[15] <= 32'h03F00FC0;
                     char22_2[16] <= 32'h03E007C0;
                     char22_2[17] <= 32'h07E007E0;
                     char22_2[18] <= 32'h07C003E0;
                     char22_2[19] <= 32'h0FC003F0;
                     char22_2[20] <= 32'h0FC003F0;
                     char22_2[21] <= 32'h0FC003F0;
                     char22_2[22] <= 32'h1F8001F8;
                     char22_2[23] <= 32'h1F8001F8;
                     char22_2[24] <= 32'h1F8001F8;
                     char22_2[25] <= 32'h1F8001F8;
                     char22_2[26] <= 32'h1F8001F8;
                     char22_2[27] <= 32'h3F8001F8;
                     char22_2[28] <= 32'h3F8001F8;
                     char22_2[29] <= 32'h3F8001F8;
                     char22_2[30] <= 32'h3F8001F8;
                     char22_2[31] <= 32'h3F8001F8;
                     char22_2[32] <= 32'h3F8001F8;
                     char22_2[33] <= 32'h3F8001F8;
                     char22_2[34] <= 32'h3F8001F8;
                     char22_2[35] <= 32'h3F8001F8;
                     char22_2[36] <= 32'h3F8001F8;
                     char22_2[37] <= 32'h1F8001F8;
                     char22_2[38] <= 32'h1F8001F8;
                     char22_2[39] <= 32'h1F8001F8;
                     char22_2[40] <= 32'h1F8001F8;
                     char22_2[41] <= 32'h1F8001F0;
                     char22_2[42] <= 32'h0F8003F0;
                     char22_2[43] <= 32'h0FC003F0;
                     char22_2[44] <= 32'h0FC003F0;
                     char22_2[45] <= 32'h07C003E0;
                     char22_2[46] <= 32'h07E007E0;
                     char22_2[47] <= 32'h03E007C0;
                     char22_2[48] <= 32'h03F00FC0;
                     char22_2[49] <= 32'h01F00F80;
                     char22_2[50] <= 32'h00F81F00;
                     char22_2[51] <= 32'h007E7E00;
                     char22_2[52] <= 32'h003FFC00;
                     char22_2[53] <= 32'h000FF000;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//0
                 4'd1: begin
                     char22_2[  0] <= 32'h00000000;
                     char22_2[  1] <= 32'h00000000;
                     char22_2[  2] <= 32'h00000000;
                     char22_2[  3] <= 32'h00000000;
                     char22_2[  4] <= 32'h00000000;
                     char22_2[  5] <= 32'h00000000;
                     char22_2[  6] <= 32'h00000000;
                     char22_2[  7] <= 32'h00000000;
                     char22_2[  8] <= 32'h00000000;
                     char22_2[  9] <= 32'h00000000;
                     char22_2[10] <= 32'h0000E000;
                     char22_2[11] <= 32'h0001E000;
                     char22_2[12] <= 32'h0003E000;
                     char22_2[13] <= 32'h001FE000;
                     char22_2[14] <= 32'h03FFE000;
                     char22_2[15] <= 32'h03FFE000;
                     char22_2[16] <= 32'h0007E000;
                     char22_2[17] <= 32'h0007E000;
                     char22_2[18] <= 32'h0007E000;
                     char22_2[19] <= 32'h0007E000;
                     char22_2[20] <= 32'h0007E000;
                     char22_2[21] <= 32'h0007E000;
                     char22_2[22] <= 32'h0007E000;
                     char22_2[23] <= 32'h0007E000;
                     char22_2[24] <= 32'h0007E000;
                     char22_2[25] <= 32'h0007E000;
                     char22_2[26] <= 32'h0007E000;
                     char22_2[27] <= 32'h0007E000;
                     char22_2[28] <= 32'h0007E000;
                     char22_2[29] <= 32'h0007E000;
                     char22_2[30] <= 32'h0007E000;
                     char22_2[31] <= 32'h0007E000;
                     char22_2[32] <= 32'h0007E000;
                     char22_2[33] <= 32'h0007E000;
                     char22_2[34] <= 32'h0007E000;
                     char22_2[35] <= 32'h0007E000;
                     char22_2[36] <= 32'h0007E000;
                     char22_2[37] <= 32'h0007E000;
                     char22_2[38] <= 32'h0007E000;
                     char22_2[39] <= 32'h0007E000;
                     char22_2[40] <= 32'h0007E000;
                     char22_2[41] <= 32'h0007E000;
                     char22_2[42] <= 32'h0007E000;
                     char22_2[43] <= 32'h0007E000;
                     char22_2[44] <= 32'h0007E000;
                     char22_2[45] <= 32'h0007E000;
                     char22_2[46] <= 32'h0007E000;
                     char22_2[47] <= 32'h0007E000;
                     char22_2[48] <= 32'h0007E000;
                     char22_2[49] <= 32'h0007E000;
                     char22_2[50] <= 32'h0007E000;
                     char22_2[51] <= 32'h000FF800;
                     char22_2[52] <= 32'h03FFFFC0;
                     char22_2[53] <= 32'h03FFFFC0;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//1
                 4'd2: begin
                     char22_2[  0] <= 32'h00000000;
                     char22_2[  1] <= 32'h00000000;
                     char22_2[  2] <= 32'h00000000;
                     char22_2[  3] <= 32'h00000000;
                     char22_2[  4] <= 32'h00000000;
                     char22_2[  5] <= 32'h00000000;
                     char22_2[  6] <= 32'h00000000;
                     char22_2[  7] <= 32'h00000000;
                     char22_2[  8] <= 32'h00000000;
                     char22_2[  9] <= 32'h00000000;
                     char22_2[10] <= 32'h001FFC00;
                     char22_2[11] <= 32'h007FFF00;
                     char22_2[12] <= 32'h01F83F80;
                     char22_2[13] <= 32'h03E00FC0;
                     char22_2[14] <= 32'h07C007E0;
                     char22_2[15] <= 32'h078007E0;
                     char22_2[16] <= 32'h0F8003F0;
                     char22_2[17] <= 32'h0F8003F0;
                     char22_2[18] <= 32'h1F8003F0;
                     char22_2[19] <= 32'h1F8003F0;
                     char22_2[20] <= 32'h1FC003F0;
                     char22_2[21] <= 32'h1FC003F0;
                     char22_2[22] <= 32'h1FC003F0;
                     char22_2[23] <= 32'h0FC003F0;
                     char22_2[24] <= 32'h07C003F0;
                     char22_2[25] <= 32'h000003E0;
                     char22_2[26] <= 32'h000007E0;
                     char22_2[27] <= 32'h000007E0;
                     char22_2[28] <= 32'h00000FC0;
                     char22_2[29] <= 32'h00000F80;
                     char22_2[30] <= 32'h00001F80;
                     char22_2[31] <= 32'h00003F00;
                     char22_2[32] <= 32'h00003E00;
                     char22_2[33] <= 32'h00007C00;
                     char22_2[34] <= 32'h0000F800;
                     char22_2[35] <= 32'h0001F000;
                     char22_2[36] <= 32'h0003E000;
                     char22_2[37] <= 32'h0007C000;
                     char22_2[38] <= 32'h000F8000;
                     char22_2[39] <= 32'h001F0000;
                     char22_2[40] <= 32'h003E0000;
                     char22_2[41] <= 32'h007C0000;
                     char22_2[42] <= 32'h00F80000;
                     char22_2[43] <= 32'h01F00038;
                     char22_2[44] <= 32'h01E00038;
                     char22_2[45] <= 32'h03C00070;
                     char22_2[46] <= 32'h07800070;
                     char22_2[47] <= 32'h0F8000F0;
                     char22_2[48] <= 32'h0F0000F0;
                     char22_2[49] <= 32'h1E0003F0;
                     char22_2[50] <= 32'h3FFFFFF0;
                     char22_2[51] <= 32'h3FFFFFF0;
                     char22_2[52] <= 32'h3FFFFFE0;
                     char22_2[53] <= 32'h3FFFFFE0;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//2
                 4'd3: begin
                     char22_2[  0] <= 32'h00000000;
                     char22_2[  1] <= 32'h00000000;
                     char22_2[  2] <= 32'h00000000;
                     char22_2[  3] <= 32'h00000000;
                     char22_2[  4] <= 32'h00000000;
                     char22_2[  5] <= 32'h00000000;
                     char22_2[  6] <= 32'h00000000;
                     char22_2[  7] <= 32'h00000000;
                     char22_2[  8] <= 32'h00000000;
                     char22_2[  9] <= 32'h00000000;
                     char22_2[10] <= 32'h003FF000;
                     char22_2[11] <= 32'h00FFFC00;
                     char22_2[12] <= 32'h01F07E00;
                     char22_2[13] <= 32'h03C03F00;
                     char22_2[14] <= 32'h07801F80;
                     char22_2[15] <= 32'h0F800FC0;
                     char22_2[16] <= 32'h0F800FC0;
                     char22_2[17] <= 32'h0F8007E0;
                     char22_2[18] <= 32'h0FC007E0;
                     char22_2[19] <= 32'h0FC007E0;
                     char22_2[20] <= 32'h0FC007E0;
                     char22_2[21] <= 32'h07C007E0;
                     char22_2[22] <= 32'h000007E0;
                     char22_2[23] <= 32'h000007E0;
                     char22_2[24] <= 32'h000007C0;
                     char22_2[25] <= 32'h00000FC0;
                     char22_2[26] <= 32'h00000F80;
                     char22_2[27] <= 32'h00001F00;
                     char22_2[28] <= 32'h00007E00;
                     char22_2[29] <= 32'h0003FC00;
                     char22_2[30] <= 32'h001FF000;
                     char22_2[31] <= 32'h001FFC00;
                     char22_2[32] <= 32'h0000FF00;
                     char22_2[33] <= 32'h00001F80;
                     char22_2[34] <= 32'h00000FC0;
                     char22_2[35] <= 32'h000007E0;
                     char22_2[36] <= 32'h000003E0;
                     char22_2[37] <= 32'h000003F0;
                     char22_2[38] <= 32'h000003F0;
                     char22_2[39] <= 32'h000001F0;
                     char22_2[40] <= 32'h000001F8;
                     char22_2[41] <= 32'h000001F8;
                     char22_2[42] <= 32'h078001F8;
                     char22_2[43] <= 32'h0FC001F8;
                     char22_2[44] <= 32'h1FC001F8;
                     char22_2[45] <= 32'h1FC003F0;
                     char22_2[46] <= 32'h1FC003F0;
                     char22_2[47] <= 32'h1FC003E0;
                     char22_2[48] <= 32'h0F8007E0;
                     char22_2[49] <= 32'h0F8007C0;
                     char22_2[50] <= 32'h07C01F80;
                     char22_2[51] <= 32'h03F07F00;
                     char22_2[52] <= 32'h01FFFE00;
                     char22_2[53] <= 32'h003FF000;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//3
                 4'd4: begin
                     char22_2[  0] <= 32'h00000000;
                     char22_2[  1] <= 32'h00000000;
                     char22_2[  2] <= 32'h00000000;
                     char22_2[  3] <= 32'h00000000;
                     char22_2[  4] <= 32'h00000000;
                     char22_2[  5] <= 32'h00000000;
                     char22_2[  6] <= 32'h00000000;
                     char22_2[  7] <= 32'h00000000;
                     char22_2[  8] <= 32'h00000000;
                     char22_2[  9] <= 32'h00000000;
                     char22_2[10] <= 32'h00001F00;
                     char22_2[11] <= 32'h00001F00;
                     char22_2[12] <= 32'h00003F00;
                     char22_2[13] <= 32'h00003F00;
                     char22_2[14] <= 32'h00007F00;
                     char22_2[15] <= 32'h0000FF00;
                     char22_2[16] <= 32'h0000FF00;
                     char22_2[17] <= 32'h0001FF00;
                     char22_2[18] <= 32'h0003FF00;
                     char22_2[19] <= 32'h0003BF00;
                     char22_2[20] <= 32'h0007BF00;
                     char22_2[21] <= 32'h00073F00;
                     char22_2[22] <= 32'h000F3F00;
                     char22_2[23] <= 32'h001E3F00;
                     char22_2[24] <= 32'h001C3F00;
                     char22_2[25] <= 32'h003C3F00;
                     char22_2[26] <= 32'h00783F00;
                     char22_2[27] <= 32'h00783F00;
                     char22_2[28] <= 32'h00F03F00;
                     char22_2[29] <= 32'h00E03F00;
                     char22_2[30] <= 32'h01E03F00;
                     char22_2[31] <= 32'h03C03F00;
                     char22_2[32] <= 32'h03803F00;
                     char22_2[33] <= 32'h07803F00;
                     char22_2[34] <= 32'h0F003F00;
                     char22_2[35] <= 32'h0F003F00;
                     char22_2[36] <= 32'h1E003F00;
                     char22_2[37] <= 32'h1C003F00;
                     char22_2[38] <= 32'h3C003F00;
                     char22_2[39] <= 32'h7FFFFFFE;
                     char22_2[40] <= 32'h7FFFFFFE;
                     char22_2[41] <= 32'h00003F00;
                     char22_2[42] <= 32'h00003F00;
                     char22_2[43] <= 32'h00003F00;
                     char22_2[44] <= 32'h00003F00;
                     char22_2[45] <= 32'h00003F00;
                     char22_2[46] <= 32'h00003F00;
                     char22_2[47] <= 32'h00003F00;
                     char22_2[48] <= 32'h00003F00;
                     char22_2[49] <= 32'h00003F00;
                     char22_2[50] <= 32'h00003F00;
                     char22_2[51] <= 32'h00007F80;
                     char22_2[52] <= 32'h000FFFFC;
                     char22_2[53] <= 32'h000FFFFC;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//4
                 4'd5: begin
                     char22_2[  0] <= 32'h00000000;
                     char22_2[  1] <= 32'h00000000;
                     char22_2[  2] <= 32'h00000000;
                     char22_2[  3] <= 32'h00000000;
                     char22_2[  4] <= 32'h00000000;
                     char22_2[  5] <= 32'h00000000;
                     char22_2[  6] <= 32'h00000000;
                     char22_2[  7] <= 32'h00000000;
                     char22_2[  8] <= 32'h00000000;
                     char22_2[  9] <= 32'h00000000;
                     char22_2[10] <= 32'h00000000;
                     char22_2[11] <= 32'h03FFFFF0;
                     char22_2[12] <= 32'h03FFFFF0;
                     char22_2[13] <= 32'h03FFFFF0;
                     char22_2[14] <= 32'h03FFFFE0;
                     char22_2[15] <= 32'h03800000;
                     char22_2[16] <= 32'h03800000;
                     char22_2[17] <= 32'h03800000;
                     char22_2[18] <= 32'h03800000;
                     char22_2[19] <= 32'h03800000;
                     char22_2[20] <= 32'h07800000;
                     char22_2[21] <= 32'h07800000;
                     char22_2[22] <= 32'h07800000;
                     char22_2[23] <= 32'h07800000;
                     char22_2[24] <= 32'h07800000;
                     char22_2[25] <= 32'h07800000;
                     char22_2[26] <= 32'h078FF800;
                     char22_2[27] <= 32'h073FFE00;
                     char22_2[28] <= 32'h077FFF80;
                     char22_2[29] <= 32'h07FC3F80;
                     char22_2[30] <= 32'h07E00FC0;
                     char22_2[31] <= 32'h07C007E0;
                     char22_2[32] <= 32'h078007E0;
                     char22_2[33] <= 32'h078003F0;
                     char22_2[34] <= 32'h000003F0;
                     char22_2[35] <= 32'h000001F0;
                     char22_2[36] <= 32'h000001F8;
                     char22_2[37] <= 32'h000001F8;
                     char22_2[38] <= 32'h000001F8;
                     char22_2[39] <= 32'h000001F8;
                     char22_2[40] <= 32'h000001F8;
                     char22_2[41] <= 32'h078001F8;
                     char22_2[42] <= 32'h0FC001F8;
                     char22_2[43] <= 32'h1FC001F0;
                     char22_2[44] <= 32'h1FC001F0;
                     char22_2[45] <= 32'h1FC003F0;
                     char22_2[46] <= 32'h1F8003F0;
                     char22_2[47] <= 32'h1F8003E0;
                     char22_2[48] <= 32'h0F8007E0;
                     char22_2[49] <= 32'h078007C0;
                     char22_2[50] <= 32'h07C01F80;
                     char22_2[51] <= 32'h03F83F00;
                     char22_2[52] <= 32'h00FFFE00;
                     char22_2[53] <= 32'h003FF800;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//5
                 4'd6: begin
                     char22_2[0] <= 32'h00000000;
                     char22_2[1] <= 32'h00000000;
                     char22_2[2] <= 32'h00000000;
                     char22_2[3] <= 32'h00000000;
                     char22_2[4] <= 32'h00000000;
                     char22_2[5] <= 32'h00000000;
                     char22_2[6] <= 32'h00000000;
                     char22_2[7] <= 32'h00000000;
                     char22_2[8] <= 32'h00000000;
                     char22_2[9] <= 32'h00000000;
                     char22_2[10] <= 32'h0007FE00;
                     char22_2[11] <= 32'h001FFF80;
                     char22_2[12] <= 32'h003F0FC0;
                     char22_2[13] <= 32'h007C07C0;
                     char22_2[14] <= 32'h00F807E0;
                     char22_2[15] <= 32'h01F007E0;
                     char22_2[16] <= 32'h03E007E0;
                     char22_2[17] <= 32'h03C007E0;
                     char22_2[18] <= 32'h07C003C0;
                     char22_2[19] <= 32'h07C00000;
                     char22_2[20] <= 32'h0FC00000;
                     char22_2[21] <= 32'h0F800000;
                     char22_2[22] <= 32'h0F800000;
                     char22_2[23] <= 32'h1F800000;
                     char22_2[24] <= 32'h1F800000;
                     char22_2[25] <= 32'h1F800000;
                     char22_2[26] <= 32'h1F87FE00;
                     char22_2[27] <= 32'h1F9FFF80;
                     char22_2[28] <= 32'h1FBFFFC0;
                     char22_2[29] <= 32'h3FFE1FC0;
                     char22_2[30] <= 32'h3FF807E0;
                     char22_2[31] <= 32'h3FE003F0;
                     char22_2[32] <= 32'h3FE003F0;
                     char22_2[33] <= 32'h3FC001F8;
                     char22_2[34] <= 32'h3F8001F8;
                     char22_2[35] <= 32'h3F8001F8;
                     char22_2[36] <= 32'h3F8000F8;
                     char22_2[37] <= 32'h3F8000F8;
                     char22_2[38] <= 32'h3F8000F8;
                     char22_2[39] <= 32'h1F8000F8;
                     char22_2[40] <= 32'h1F8000F8;
                     char22_2[41] <= 32'h1F8000F8;
                     char22_2[42] <= 32'h1F8000F8;
                     char22_2[43] <= 32'h1F8000F8;
                     char22_2[44] <= 32'h0FC001F8;
                     char22_2[45] <= 32'h0FC001F8;
                     char22_2[46] <= 32'h0FC001F0;
                     char22_2[47] <= 32'h07E001F0;
                     char22_2[48] <= 32'h03E003E0;
                     char22_2[49] <= 32'h03F003E0;
                     char22_2[50] <= 32'h01F807C0;
                     char22_2[51] <= 32'h00FE1F80;
                     char22_2[52] <= 32'h007FFE00;
                     char22_2[53] <= 32'h001FF800;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//6
                 4'd7: begin
                     char22_2[0] <= 32'h00000000;
                     char22_2[1] <= 32'h00000000;
                     char22_2[2] <= 32'h00000000;
                     char22_2[3] <= 32'h00000000;
                     char22_2[4] <= 32'h00000000;
                     char22_2[5] <= 32'h00000000;
                     char22_2[6] <= 32'h00000000;
                     char22_2[7] <= 32'h00000000;
                     char22_2[8] <= 32'h00000000;
                     char22_2[9] <= 32'h00000000;
                     char22_2[10] <= 32'h00000000;
                     char22_2[11] <= 32'h07FFFFF8;
                     char22_2[12] <= 32'h07FFFFF8;
                     char22_2[13] <= 32'h07FFFFF8;
                     char22_2[14] <= 32'h0FFFFFF0;
                     char22_2[15] <= 32'h0FC000E0;
                     char22_2[16] <= 32'h0F8001E0;
                     char22_2[17] <= 32'h0F0001C0;
                     char22_2[18] <= 32'h0E0003C0;
                     char22_2[19] <= 32'h0E000780;
                     char22_2[20] <= 32'h1E000780;
                     char22_2[21] <= 32'h1C000F00;
                     char22_2[22] <= 32'h00000F00;
                     char22_2[23] <= 32'h00001E00;
                     char22_2[24] <= 32'h00001E00;
                     char22_2[25] <= 32'h00003C00;
                     char22_2[26] <= 32'h00003C00;
                     char22_2[27] <= 32'h00007800;
                     char22_2[28] <= 32'h00007800;
                     char22_2[29] <= 32'h0000F800;
                     char22_2[30] <= 32'h0000F000;
                     char22_2[31] <= 32'h0001F000;
                     char22_2[32] <= 32'h0001E000;
                     char22_2[33] <= 32'h0003E000;
                     char22_2[34] <= 32'h0003E000;
                     char22_2[35] <= 32'h0003E000;
                     char22_2[36] <= 32'h0007C000;
                     char22_2[37] <= 32'h0007C000;
                     char22_2[38] <= 32'h0007C000;
                     char22_2[39] <= 32'h000FC000;
                     char22_2[40] <= 32'h000FC000;
                     char22_2[41] <= 32'h000FC000;
                     char22_2[42] <= 32'h000FC000;
                     char22_2[43] <= 32'h001FC000;
                     char22_2[44] <= 32'h001FC000;
                     char22_2[45] <= 32'h001FC000;
                     char22_2[46] <= 32'h001FC000;
                     char22_2[47] <= 32'h001FC000;
                     char22_2[48] <= 32'h001FC000;
                     char22_2[49] <= 32'h001FC000;
                     char22_2[50] <= 32'h001FC000;
                     char22_2[51] <= 32'h001FC000;
                     char22_2[52] <= 32'h001FC000;
                     char22_2[53] <= 32'h000F8000;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//7
                 4'd8: begin
                     char22_2[0] <= 32'h00000000;
                     char22_2[1] <= 32'h00000000;
                     char22_2[2] <= 32'h00000000;
                     char22_2[3] <= 32'h00000000;
                     char22_2[4] <= 32'h00000000;
                     char22_2[5] <= 32'h00000000;
                     char22_2[6] <= 32'h00000000;
                     char22_2[7] <= 32'h00000000;
                     char22_2[8] <= 32'h00000000;
                     char22_2[9] <= 32'h00000000;
                     char22_2[10] <= 32'h003FF800;
                     char22_2[11] <= 32'h00FFFE00;
                     char22_2[12] <= 32'h01F81F80;
                     char22_2[13] <= 32'h03E00FC0;
                     char22_2[14] <= 32'h07C003E0;
                     char22_2[15] <= 32'h0F8003E0;
                     char22_2[16] <= 32'h0F8001F0;
                     char22_2[17] <= 32'h1F0001F0;
                     char22_2[18] <= 32'h1F0001F0;
                     char22_2[19] <= 32'h1F0001F0;
                     char22_2[20] <= 32'h1F0001F0;
                     char22_2[21] <= 32'h1F0001F0;
                     char22_2[22] <= 32'h1F8001F0;
                     char22_2[23] <= 32'h1FC001F0;
                     char22_2[24] <= 32'h0FC001F0;
                     char22_2[25] <= 32'h0FF003E0;
                     char22_2[26] <= 32'h07F803C0;
                     char22_2[27] <= 32'h03FE0F80;
                     char22_2[28] <= 32'h01FF9F00;
                     char22_2[29] <= 32'h00FFFE00;
                     char22_2[30] <= 32'h003FF800;
                     char22_2[31] <= 32'h007FFC00;
                     char22_2[32] <= 32'h01F7FF00;
                     char22_2[33] <= 32'h03E1FF80;
                     char22_2[34] <= 32'h07C07FC0;
                     char22_2[35] <= 32'h0F801FE0;
                     char22_2[36] <= 32'h0F800FE0;
                     char22_2[37] <= 32'h1F0007F0;
                     char22_2[38] <= 32'h1F0003F0;
                     char22_2[39] <= 32'h3E0001F8;
                     char22_2[40] <= 32'h3E0001F8;
                     char22_2[41] <= 32'h3E0001F8;
                     char22_2[42] <= 32'h3E0000F8;
                     char22_2[43] <= 32'h3E0000F8;
                     char22_2[44] <= 32'h3E0000F8;
                     char22_2[45] <= 32'h3E0000F8;
                     char22_2[46] <= 32'h1F0001F0;
                     char22_2[47] <= 32'h1F0001F0;
                     char22_2[48] <= 32'h0F8003E0;
                     char22_2[49] <= 32'h0FC003E0;
                     char22_2[50] <= 32'h07E007C0;
                     char22_2[51] <= 32'h01F83F80;
                     char22_2[52] <= 32'h00FFFE00;
                     char22_2[53] <= 32'h003FF800;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//8
                 4'd9: begin
                     char22_2[0] <= 32'h00000000;
                     char22_2[1] <= 32'h00000000;
                     char22_2[2] <= 32'h00000000;
                     char22_2[3] <= 32'h00000000;
                     char22_2[4] <= 32'h00000000;
                     char22_2[5] <= 32'h00000000;
                     char22_2[6] <= 32'h00000000;
                     char22_2[7] <= 32'h00000000;
                     char22_2[8] <= 32'h00000000;
                     char22_2[9] <= 32'h00000000;
                     char22_2[10] <= 32'h003FF000;
                     char22_2[11] <= 32'h00FFFC00;
                     char22_2[12] <= 32'h01F83F00;
                     char22_2[13] <= 32'h03E01F80;
                     char22_2[14] <= 32'h07C00F80;
                     char22_2[15] <= 32'h0FC007C0;
                     char22_2[16] <= 32'h0F8003E0;
                     char22_2[17] <= 32'h1F8003E0;
                     char22_2[18] <= 32'h1F0003F0;
                     char22_2[19] <= 32'h1F0003F0;
                     char22_2[20] <= 32'h3F0001F0;
                     char22_2[21] <= 32'h3F0001F0;
                     char22_2[22] <= 32'h3F0001F8;
                     char22_2[23] <= 32'h3F0001F8;
                     char22_2[24] <= 32'h3F0001F8;
                     char22_2[25] <= 32'h3F0001F8;
                     char22_2[26] <= 32'h3F0001F8;
                     char22_2[27] <= 32'h3F0001F8;
                     char22_2[28] <= 32'h3F0003F8;
                     char22_2[29] <= 32'h1F8003F8;
                     char22_2[30] <= 32'h1F8007F8;
                     char22_2[31] <= 32'h1F800FF8;
                     char22_2[32] <= 32'h0FC01FF8;
                     char22_2[33] <= 32'h0FE03FF8;
                     char22_2[34] <= 32'h07F8FDF8;
                     char22_2[35] <= 32'h03FFF9F8;
                     char22_2[36] <= 32'h01FFF1F8;
                     char22_2[37] <= 32'h003F83F8;
                     char22_2[38] <= 32'h000003F0;
                     char22_2[39] <= 32'h000003F0;
                     char22_2[40] <= 32'h000003F0;
                     char22_2[41] <= 32'h000003F0;
                     char22_2[42] <= 32'h000007E0;
                     char22_2[43] <= 32'h000007E0;
                     char22_2[44] <= 32'h000007C0;
                     char22_2[45] <= 32'h03C007C0;
                     char22_2[46] <= 32'h07C00F80;
                     char22_2[47] <= 32'h0FE00F80;
                     char22_2[48] <= 32'h0FE01F00;
                     char22_2[49] <= 32'h0FE03E00;
                     char22_2[50] <= 32'h07E07E00;
                     char22_2[51] <= 32'h07F1F800;
                     char22_2[52] <= 32'h03FFF000;
                     char22_2[53] <= 32'h00FFC000;
                     char22_2[54] <= 32'h00000000;
                     char22_2[55] <= 32'h00000000;
                     char22_2[56] <= 32'h00000000;
                     char22_2[57] <= 32'h00000000;
                     char22_2[58] <= 32'h00000000;
                     char22_2[59] <= 32'h00000000;
                     char22_2[60] <= 32'h00000000;
                     char22_2[61] <= 32'h00000000;
                     char22_2[62] <= 32'h00000000;
                     char22_2[63] <= 32'h00000000;
                 end//9
                 default: begin
                     char22_2[0] <= char22_2[0];
                     char22_2[1] <= char22_2[1];
                     char22_2[2] <= char22_2[2];
                     char22_2[3] <= char22_2[3];
                     char22_2[4] <= char22_2[4];
                     char22_2[5] <= char22_2[5];
                     char22_2[6] <= char22_2[6];
                     char22_2[7] <= char22_2[7];
                     char22_2[8] <= char22_2[8];
                     char22_2[9] <= char22_2[9];
                     char22_2[10] <= char22_2[10];
                     char22_2[11] <= char22_2[11];
                     char22_2[12] <= char22_2[12];
                     char22_2[13] <= char22_2[13];
                     char22_2[14] <= char22_2[14];
                     char22_2[15] <= char22_2[15];
                     char22_2[16] <= char22_2[16];
                     char22_2[17] <= char22_2[17];
                     char22_2[18] <= char22_2[18];
                     char22_2[19] <= char22_2[19];
                     char22_2[20] <= char22_2[20];
                     char22_2[21] <= char22_2[21];
                     char22_2[22] <= char22_2[22];
                     char22_2[23] <= char22_2[23];
                     char22_2[24] <= char22_2[24];
                     char22_2[25] <= char22_2[25];
                     char22_2[26] <= char22_2[26];
                     char22_2[27] <= char22_2[27];
                     char22_2[28] <= char22_2[28];
                     char22_2[29] <= char22_2[29];
                     char22_2[30] <= char22_2[30];
                     char22_2[31] <= char22_2[31];
                     char22_2[32] <= char22_2[32];
                     char22_2[33] <= char22_2[33];
                     char22_2[34] <= char22_2[34];
                     char22_2[35] <= char22_2[35];
                     char22_2[36] <= char22_2[36];
                     char22_2[37] <= char22_2[37];
                     char22_2[38] <= char22_2[38];
                     char22_2[39] <= char22_2[39];
                     char22_2[40] <= char22_2[40];
                     char22_2[41] <= char22_2[41];
                     char22_2[42] <= char22_2[42];
                     char22_2[43] <= char22_2[43];
                     char22_2[44] <= char22_2[44];
                     char22_2[45] <= char22_2[45];
                     char22_2[46] <= char22_2[46];
                     char22_2[47] <= char22_2[47];
                     char22_2[48] <= char22_2[48];
                     char22_2[49] <= char22_2[49];
                     char22_2[50] <= char22_2[50];
                     char22_2[51] <= char22_2[51];
                     char22_2[52] <= char22_2[52];
                     char22_2[53] <= char22_2[53];
                     char22_2[54] <= char22_2[54];
                     char22_2[55] <= char22_2[55];
                     char22_2[56] <= char22_2[56];
                     char22_2[57] <= char22_2[57];
                     char22_2[58] <= char22_2[58];
                     char22_2[59] <= char22_2[59];
                     char22_2[60] <= char22_2[60];
                     char22_2[61] <= char22_2[61];
                     char22_2[62] <= char22_2[62];
                     char22_2[63] <= char22_2[63];
                 end
             endcase
     
    
         case((li - onekm*(li/onekm))/diankm)
                    4'd0: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h000FF000000000000000000000000000;
                          char22_4[11] <= 128'h003FFC00000000000000000000000000;
                          char22_4[12] <= 128'h007E7E00800000000000000000000000;
                          char22_4[13] <= 128'h00F81F00000000000000000000000000;
                          char22_4[14] <= 128'h01F00F80000000000000000000000000;
                          char22_4[15] <= 128'h03F00FC0000000000000000000000000;
                          char22_4[16] <= 128'h03E007C0000000000000000000000000;
                          char22_4[17] <= 128'h07E007E0000000000000000000000000;
                          char22_4[18] <= 128'h07C003E0000000000000000000000000;
                          char22_4[19] <= 128'h0FC003F0000000000000000000000000;
                          char22_4[20] <= 128'h0FC003F0000000000000000000000000;
                          char22_4[21] <= 128'h0FC003F0000000000000000000000000;
                          char22_4[22] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[23] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[24] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[25] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[26] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[27] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[28] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[29] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[30] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[31] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[32] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[33] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[34] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[35] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[36] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[37] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[38] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[39] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[40] <= 128'h1F8001F8000000000000000000000000;
                          char22_4[41] <= 128'h1F8001F0000000000000000000000000;
                          char22_4[42] <= 128'h0F8003F0000000000000000000000000;
                          char22_4[43] <= 128'h0FC003F0000000000000000000000000;
                          char22_4[44] <= 128'h0FC003F0000000000000000000000000;
                          char22_4[45] <= 128'h07C003E0000000000000000000000000;
                          char22_4[46] <= 128'h07E007E0000000000000000000000000;
                          char22_4[47] <= 128'h03E007C0000000000000000000000000;
                          char22_4[48] <= 128'h03F00FC0000000000000000000000000;
                          char22_4[49] <= 128'h01F00F80000000000000000000000000;
                          char22_4[50] <= 128'h00F81F00000000000000000000000000;
                          char22_4[51] <= 128'h007E7E00000000000000000000000000;
                          char22_4[52] <= 128'h003FFC00000000000000000000000000;
                          char22_4[53] <= 128'h000FF000000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//0
                    4'd1: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h0000E000000000000000000000000000;
                          char22_4[11] <= 128'h0001E000000000000000000000000000;
                          char22_4[12] <= 128'h0003E000000000000000000000000000;
                          char22_4[13] <= 128'h001FE000000000000000000000000000;
                          char22_4[14] <= 128'h03FFE000000000000000000000000000;
                          char22_4[15] <= 128'h03FFE000000000000000000000000000;
                          char22_4[16] <= 128'h0007E000000000000000000000000000;
                          char22_4[17] <= 128'h0007E000000000000000000000000000;
                          char22_4[18] <= 128'h0007E000000000000000000000000000;
                          char22_4[19] <= 128'h0007E000000000000000000000000000;
                          char22_4[20] <= 128'h0007E000000000000000000000000000;
                          char22_4[21] <= 128'h0007E000000000000000000000000000;
                          char22_4[22] <= 128'h0007E000000000000000000000000000;
                          char22_4[23] <= 128'h0007E000000000000000000000000000;
                          char22_4[24] <= 128'h0007E000000000000000000000000000;
                          char22_4[25] <= 128'h0007E000000000000000000000000000;
                          char22_4[26] <= 128'h0007E000000000000000000000000000;
                          char22_4[27] <= 128'h0007E000000000000000000000000000;
                          char22_4[28] <= 128'h0007E000000000000000000000000000;
                          char22_4[29] <= 128'h0007E000000000000000000000000000;
                          char22_4[30] <= 128'h0007E000000000000000000000000000;
                          char22_4[31] <= 128'h0007E000000000000000000000000000;
                          char22_4[32] <= 128'h0007E000000000000000000000000000;
                          char22_4[33] <= 128'h0007E000000000000000000000000000;
                          char22_4[34] <= 128'h0007E000000000000000000000000000;
                          char22_4[35] <= 128'h0007E000000000000000000000000000;
                          char22_4[36] <= 128'h0007E000000000000000000000000000;
                          char22_4[37] <= 128'h0007E000000000000000000000000000;
                          char22_4[38] <= 128'h0007E000000000000000000000000000;
                          char22_4[39] <= 128'h0007E000000000000000000000000000;
                          char22_4[40] <= 128'h0007E000000000000000000000000000;
                          char22_4[41] <= 128'h0007E000000000000000000000000000;
                          char22_4[42] <= 128'h0007E000000000000000000000000000;
                          char22_4[43] <= 128'h0007E000000000000000000000000000;
                          char22_4[44] <= 128'h0007E000000000000000000000000000;
                          char22_4[45] <= 128'h0007E000000000000000000000000000;
                          char22_4[46] <= 128'h0007E000000000000000000000000000;
                          char22_4[47] <= 128'h0007E000000000000000000000000000;
                          char22_4[48] <= 128'h0007E000000000000000000000000000;
                          char22_4[49] <= 128'h0007E000000000000000000000000000;
                          char22_4[50] <= 128'h0007E000000000000000000000000000;
                          char22_4[51] <= 128'h000FF800000000000000000000000000;
                          char22_4[52] <= 128'h03FFFFC0000000000000000000000000;
                          char22_4[53] <= 128'h03FFFFC0000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//1
                    4'd2: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h001FFC00000000000000000000000000;
                          char22_4[11] <= 128'h007FFF00000000000000000000000000;
                          char22_4[12] <= 128'h01F83F80000000000000000000000000;
                          char22_4[13] <= 128'h03E00FC0000000000000000000000000;
                          char22_4[14] <= 128'h07C007E0000000000000000000000000;
                          char22_4[15] <= 128'h078007E0000000000000000000000000;
                          char22_4[16] <= 128'h0F8003F0000000000000000000000000;
                          char22_4[17] <= 128'h0F8003F0000000000000000000000000;
                          char22_4[18] <= 128'h1F8003F0000000000000000000000000;
                          char22_4[19] <= 128'h1F8003F0000000000000000000000000;
                          char22_4[20] <= 128'h1FC003F0000000000000000000000000;
                          char22_4[21] <= 128'h1FC003F0000000000000000000000000;
                          char22_4[22] <= 128'h1FC003F0000000000000000000000000;
                          char22_4[23] <= 128'h0FC003F0000000000000000000000000;
                          char22_4[24] <= 128'h07C003F0000000000000000000000000;
                          char22_4[25] <= 128'h000003E0000000000000000000000000;
                          char22_4[26] <= 128'h000007E0000000000000000000000000;
                          char22_4[27] <= 128'h000007E0000000000000000000000000;
                          char22_4[28] <= 128'h00000FC0000000000000000000000000;
                          char22_4[29] <= 128'h00000F80000000000000000000000000;
                          char22_4[30] <= 128'h00001F80000000000000000000000000;
                          char22_4[31] <= 128'h00003F00000000000000000000000000;
                          char22_4[32] <= 128'h00003E00000000000000000000000000;
                          char22_4[33] <= 128'h00007C00000000000000000000000000;
                          char22_4[34] <= 128'h0000F800000000000000000000000000;
                          char22_4[35] <= 128'h0001F000000000000000000000000000;
                          char22_4[36] <= 128'h0003E000000000000000000000000000;
                          char22_4[37] <= 128'h0007C000000000000000000000000000;
                          char22_4[38] <= 128'h000F8000000000000000000000000000;
                          char22_4[39] <= 128'h001F0000000000000000000000000000;
                          char22_4[40] <= 128'h003E0000000000000000000000000000;
                          char22_4[41] <= 128'h007C0000000000000000000000000000;
                          char22_4[42] <= 128'h00F80000000000000000000000000000;
                          char22_4[43] <= 128'h01F00038000000000000000000000000;
                          char22_4[44] <= 128'h01E00038000000000000000000000000;
                          char22_4[45] <= 128'h03C00070000000000000000000000000;
                          char22_4[46] <= 128'h07800070000000000000000000000000;
                          char22_4[47] <= 128'h0F8000F0000000000000000000000000;
                          char22_4[48] <= 128'h0F0000F0000000000000000000000000;
                          char22_4[49] <= 128'h1E0003F0000000000000000000000000;
                          char22_4[50] <= 128'h3FFFFFF0000000000000000000000000;
                          char22_4[51] <= 128'h3FFFFFF0000000000000000000000000;
                          char22_4[52] <= 128'h3FFFFFE0000000000000000000000000;
                          char22_4[53] <= 128'h3FFFFFE0000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//2
                    4'd3: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h003FF000000000000000000000000000;
                          char22_4[11] <= 128'h00FFFC00000000000000000000000000;
                          char22_4[12] <= 128'h01F07E00000000000000000000000000;
                          char22_4[13] <= 128'h03C03F00000000000000000000000000;
                          char22_4[14] <= 128'h07801F80000000000000000000000000;
                          char22_4[15] <= 128'h0F800FC0000000000000000000000000;
                          char22_4[16] <= 128'h0F800FC0000000000000000000000000;
                          char22_4[17] <= 128'h0F8007E0000000000000000000000000;
                          char22_4[18] <= 128'h0FC007E0000000000000000000000000;
                          char22_4[19] <= 128'h0FC007E0000000000000000000000000;
                          char22_4[20] <= 128'h0FC007E0000000000000000000000000;
                          char22_4[21] <= 128'h07C007E0000000000000000000000000;
                          char22_4[22] <= 128'h000007E0000000000000000000000000;
                          char22_4[23] <= 128'h000007E0000000000000000000000000;
                          char22_4[24] <= 128'h000007C0000000000000000000000000;
                          char22_4[25] <= 128'h00000FC0000000000000000000000000;
                          char22_4[26] <= 128'h00000F80000000000000000000000000;
                          char22_4[27] <= 128'h00001F00000000000000000000000000;
                          char22_4[28] <= 128'h00007E00000000000000000000000000;
                          char22_4[29] <= 128'h0003FC00000000000000000000000000;
                          char22_4[30] <= 128'h001FF000000000000000000000000000;
                          char22_4[31] <= 128'h001FFC00000000000000000000000000;
                          char22_4[32] <= 128'h0000FF00000000000000000000000000;
                          char22_4[33] <= 128'h00001F80000000000000000000000000;
                          char22_4[34] <= 128'h00000FC0000000000000000000000000;
                          char22_4[35] <= 128'h000007E0000000000000000000000000;
                          char22_4[36] <= 128'h000003E0000000000000000000000000;
                          char22_4[37] <= 128'h000003F0000000000000000000000000;
                          char22_4[38] <= 128'h000003F0000000000000000000000000;
                          char22_4[39] <= 128'h000001F0000000000000000000000000;
                          char22_4[40] <= 128'h000001F8000000000000000000000000;
                          char22_4[41] <= 128'h000001F8000000000000000000000000;
                          char22_4[42] <= 128'h078001F8000000000000000000000000;
                          char22_4[43] <= 128'h0FC001F8000000000000000000000000;
                          char22_4[44] <= 128'h1FC001F8000000000000000000000000;
                          char22_4[45] <= 128'h1FC003F0000000000000000000000000;
                          char22_4[46] <= 128'h1FC003F0000000000000000000000000;
                          char22_4[47] <= 128'h1FC003E0000000000000000000000000;
                          char22_4[48] <= 128'h0F8007E0000000000000000000000000;
                          char22_4[49] <= 128'h0F8007C0000000000000000000000000;
                          char22_4[50] <= 128'h07C01F80000000000000000000000000;
                          char22_4[51] <= 128'h03F07F00000000000000000000000000;
                          char22_4[52] <= 128'h01FFFE00000000000000000000000000;
                          char22_4[53] <= 128'h003FF000000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//3
                    4'd4: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h00001F00000000000000000000000000;
                          char22_4[11] <= 128'h00001F00000000000000000000000000;
                          char22_4[12] <= 128'h00003F00000000000000000000000000;
                          char22_4[13] <= 128'h00003F00000000000000000000000000;
                          char22_4[14] <= 128'h00007F00000000000000000000000000;
                          char22_4[15] <= 128'h0000FF00000000000000000000000000;
                          char22_4[16] <= 128'h0000FF00000000000000000000000000;
                          char22_4[17] <= 128'h0001FF00000000000000000000000000;
                          char22_4[18] <= 128'h0003FF00000000000000000000000000;
                          char22_4[19] <= 128'h0003BF00000000000000000000000000;
                          char22_4[20] <= 128'h0007BF00000000000000000000000000;
                          char22_4[21] <= 128'h00073F00000000000000000000000000;
                          char22_4[22] <= 128'h000F3F00000000000000000000000000;
                          char22_4[23] <= 128'h001E3F00000000000000000000000000;
                          char22_4[24] <= 128'h001C3F00000000000000000000000000;
                          char22_4[25] <= 128'h003C3F00000000000000000000000000;
                          char22_4[26] <= 128'h00783F00000000000000000000000000;
                          char22_4[27] <= 128'h00783F00000000000000000000000000;
                          char22_4[28] <= 128'h00F03F00000000000000000000000000;
                          char22_4[29] <= 128'h00E03F00000000000000000000000000;
                          char22_4[30] <= 128'h01E03F00000000000000000000000000;
                          char22_4[31] <= 128'h03C03F00000000000000000000000000;
                          char22_4[32] <= 128'h03803F00000000000000000000000000;
                          char22_4[33] <= 128'h07803F00000000000000000000000000;
                          char22_4[34] <= 128'h0F003F00000000000000000000000000;
                          char22_4[35] <= 128'h0F003F00000000000000000000000000;
                          char22_4[36] <= 128'h1E003F00000000000000000000000000;
                          char22_4[37] <= 128'h1C003F00000000000000000000000000;
                          char22_4[38] <= 128'h3C003F00000000000000000000000000;
                          char22_4[39] <= 128'h7FFFFFFE000000000000000000000000;
                          char22_4[40] <= 128'h7FFFFFFE000000000000000000000000;
                          char22_4[41] <= 128'h00003F00000000000000000000000000;
                          char22_4[42] <= 128'h00003F00000000000000000000000000;
                          char22_4[43] <= 128'h00003F00000000000000000000000000;
                          char22_4[44] <= 128'h00003F00000000000000000000000000;
                          char22_4[45] <= 128'h00003F00000000000000000000000000;
                          char22_4[46] <= 128'h00003F00000000000000000000000000;
                          char22_4[47] <= 128'h00003F00000000000000000000000000;
                          char22_4[48] <= 128'h00003F00000000000000000000000000;
                          char22_4[49] <= 128'h00003F00000000000000000000000000;
                          char22_4[50] <= 128'h00003F00000000000000000000000000;
                          char22_4[51] <= 128'h00007F80000000000000000000000000;
                          char22_4[52] <= 128'h000FFFFC000000000000000000000000;
                          char22_4[53] <= 128'h000FFFFC000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//4
                    4'd5: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h00000000000000000000000000000000;
                          char22_4[11] <= 128'h03FFFFF0000000000000000000000000;
                          char22_4[12] <= 128'h03FFFFF0000000000000000000000000;
                          char22_4[13] <= 128'h03FFFFF0000000000000000000000000;
                          char22_4[14] <= 128'h03FFFFE0000000000000000000000000;
                          char22_4[15] <= 128'h03800000000000000000000000000000;
                          char22_4[16] <= 128'h03800000000000000000000000000000;
                          char22_4[17] <= 128'h03800000000000000000000000000000;
                          char22_4[18] <= 128'h03800000000000000000000000000000;
                          char22_4[19] <= 128'h03800000000000000000000000000000;
                          char22_4[20] <= 128'h07800000000000000000000000000000;
                          char22_4[21] <= 128'h07800000000000000000000000000000;
                          char22_4[22] <= 128'h07800000000000000000000000000000;
                          char22_4[23] <= 128'h07800000000000000000000000000000;
                          char22_4[24] <= 128'h07800000000000000000000000000000;
                          char22_4[25] <= 128'h07800000000000000000000000000000;
                          char22_4[26] <= 128'h078FF800000000000000000000000000;
                          char22_4[27] <= 128'h073FFE00000000000000000000000000;
                          char22_4[28] <= 128'h077FFF80000000000000000000000000;
                          char22_4[29] <= 128'h07FC3F80000000000000000000000000;
                          char22_4[30] <= 128'h07E00FC0000000000000000000000000;
                          char22_4[31] <= 128'h07C007E0000000000000000000000000;
                          char22_4[32] <= 128'h078007E0000000000000000000000000;
                          char22_4[33] <= 128'h078003F0000000000000000000000000;
                          char22_4[34] <= 128'h000003F0000000000000000000000000;
                          char22_4[35] <= 128'h000001F0000000000000000000000000;
                          char22_4[36] <= 128'h000001F8000000000000000000000000;
                          char22_4[37] <= 128'h000001F8000000000000000000000000;
                          char22_4[38] <= 128'h000001F8000000000000000000000000;
                          char22_4[39] <= 128'h000001F8000000000000000000000000;
                          char22_4[40] <= 128'h000001F8000000000000000000000000;
                          char22_4[41] <= 128'h078001F8000000000000000000000000;
                          char22_4[42] <= 128'h0FC001F8000000000000000000000000;
                          char22_4[43] <= 128'h1FC001F0000000000000000000000000;
                          char22_4[44] <= 128'h1FC001F0000000000000000000000000;
                          char22_4[45] <= 128'h1FC003F0000000000000000000000000;
                          char22_4[46] <= 128'h1F8003F0000000000000000000000000;
                          char22_4[47] <= 128'h1F8003E0000000000000000000000000;
                          char22_4[48] <= 128'h0F8007E0000000000000000000000000;
                          char22_4[49] <= 128'h078007C0000000000000000000000000;
                          char22_4[50] <= 128'h07C01F80000000000000000000000000;
                          char22_4[51] <= 128'h03F83F00000000000000000000000000;
                          char22_4[52] <= 128'h00FFFE00000000000000000000000000;
                          char22_4[53] <= 128'h003FF800000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//5
                    4'd6: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h0007FE00000000000000000000000000;
                          char22_4[11] <= 128'h001FFF80000000000000000000000000;
                          char22_4[12] <= 128'h003F0FC0000000000000000000000000;
                          char22_4[13] <= 128'h007C07C0000000000000000000000000;
                          char22_4[14] <= 128'h00F807E0000000000000000000000000;
                          char22_4[15] <= 128'h01F007E0000000000000000000000000;
                          char22_4[16] <= 128'h03E007E0000000000000000000000000;
                          char22_4[17] <= 128'h03C007E0000000000000000000000000;
                          char22_4[18] <= 128'h07C003C0000000000000000000000000;
                          char22_4[19] <= 128'h07C00000000000000000000000000000;
                          char22_4[20] <= 128'h0FC00000000000000000000000000000;
                          char22_4[21] <= 128'h0F800000000000000000000000000000;
                          char22_4[22] <= 128'h0F800000000000000000000000000000;
                          char22_4[23] <= 128'h1F800000000000000000000000000000;
                          char22_4[24] <= 128'h1F800000000000000000000000000000;
                          char22_4[25] <= 128'h1F800000000000000000000000000000;
                          char22_4[26] <= 128'h1F87FE00000000000000000000000000;
                          char22_4[27] <= 128'h1F9FFF80000000000000000000000000;
                          char22_4[28] <= 128'h1FBFFFC0000000000000000000000000;
                          char22_4[29] <= 128'h3FFE1FC0000000000000000000000000;
                          char22_4[30] <= 128'h3FF807E0000000000000000000000000;
                          char22_4[31] <= 128'h3FE003F0000000000000000000000000;
                          char22_4[32] <= 128'h3FE003F0000000000000000000000000;
                          char22_4[33] <= 128'h3FC001F8000000000000000000000000;
                          char22_4[34] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[35] <= 128'h3F8001F8000000000000000000000000;
                          char22_4[36] <= 128'h3F8000F8000000000000000000000000;
                          char22_4[37] <= 128'h3F8000F8000000000000000000000000;
                          char22_4[38] <= 128'h3F8000F8000000000000000000000000;
                          char22_4[39] <= 128'h1F8000F8000000000000000000000000;
                          char22_4[40] <= 128'h1F8000F8000000000000000000000000;
                          char22_4[41] <= 128'h1F8000F8000000000000000000000000;
                          char22_4[42] <= 128'h1F8000F8000000000000000000000000;
                          char22_4[43] <= 128'h1F8000F8000000000000000000000000;
                          char22_4[44] <= 128'h0FC001F8000000000000000000000000;
                          char22_4[45] <= 128'h0FC001F8000000000000000000000000;
                          char22_4[46] <= 128'h0FC001F0000000000000000000000000;
                          char22_4[47] <= 128'h07E001F0000000000000000000000000;
                          char22_4[48] <= 128'h03E003E0000000000000000000000000;
                          char22_4[49] <= 128'h03F003E0000000000000000000000000;
                          char22_4[50] <= 128'h01F807C0000000000000000000000000;
                          char22_4[51] <= 128'h00FE1F80000000000000000000000000;
                          char22_4[52] <= 128'h007FFE00000000000000000000000000;
                          char22_4[53] <= 128'h001FF800000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//6
                    4'd7: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h00000000000000000000000000000000;
                          char22_4[11] <= 128'h07FFFFF8000000000000000000000000;
                          char22_4[12] <= 128'h07FFFFF8000000000000000000000000;
                          char22_4[13] <= 128'h07FFFFF8000000000000000000000000;
                          char22_4[14] <= 128'h0FFFFFF0000000000000000000000000;
                          char22_4[15] <= 128'h0FC000E0000000000000000000000000;
                          char22_4[16] <= 128'h0F8001E0000000000000000000000000;
                          char22_4[17] <= 128'h0F0001C0000000000000000000000000;
                          char22_4[18] <= 128'h0E0003C0000000000000000000000000;
                          char22_4[19] <= 128'h0E000780000000000000000000000000;
                          char22_4[20] <= 128'h1E000780000000000000000000000000;
                          char22_4[21] <= 128'h1C000F00000000000000000000000000;
                          char22_4[22] <= 128'h00000F00000000000000000000000000;
                          char22_4[23] <= 128'h00001E00000000000000000000000000;
                          char22_4[24] <= 128'h00001E00000000000000000000000000;
                          char22_4[25] <= 128'h00003C00000000000000000000000000;
                          char22_4[26] <= 128'h00003C00000000000000000000000000;
                          char22_4[27] <= 128'h00007800000000000000000000000000;
                          char22_4[28] <= 128'h00007800000000000000000000000000;
                          char22_4[29] <= 128'h0000F800000000000000000000000000;
                          char22_4[30] <= 128'h0000F000000000000000000000000000;
                          char22_4[31] <= 128'h0001F000000000000000000000000000;
                          char22_4[32] <= 128'h0001E000000000000000000000000000;
                          char22_4[33] <= 128'h0003E000000000000000000000000000;
                          char22_4[34] <= 128'h0003E000000000000000000000000000;
                          char22_4[35] <= 128'h0003E000000000000000000000000000;
                          char22_4[36] <= 128'h0007C000000000000000000000000000;
                          char22_4[37] <= 128'h0007C000000000000000000000000000;
                          char22_4[38] <= 128'h0007C000000000000000000000000000;
                          char22_4[39] <= 128'h000FC000000000000000000000000000;
                          char22_4[40] <= 128'h000FC000000000000000000000000000;
                          char22_4[41] <= 128'h000FC000000000000000000000000000;
                          char22_4[42] <= 128'h000FC000000000000000000000000000;
                          char22_4[43] <= 128'h001FC000000000000000000000000000;
                          char22_4[44] <= 128'h001FC000000000000000000000000000;
                          char22_4[45] <= 128'h001FC000000000000000000000000000;
                          char22_4[46] <= 128'h001FC000000000000000000000000000;
                          char22_4[47] <= 128'h001FC000000000000000000000000000;
                          char22_4[48] <= 128'h001FC000000000000000000000000000;
                          char22_4[49] <= 128'h001FC000000000000000000000000000;
                          char22_4[50] <= 128'h001FC000000000000000000000000000;
                          char22_4[51] <= 128'h001FC000000000000000000000000000;
                          char22_4[52] <= 128'h001FC000000000000000000000000000;
                          char22_4[53] <= 128'h000F8000000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//7
                    4'd8: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h003FF800000000000000000000000000;
                          char22_4[11] <= 128'h00FFFE00000000000000000000000000;
                          char22_4[12] <= 128'h01F81F80000000000000000000000000;
                          char22_4[13] <= 128'h03E00FC0000000000000000000000000;
                          char22_4[14] <= 128'h07C003E0000000000000000000000000;
                          char22_4[15] <= 128'h0F8003E0000000000000000000000000;
                          char22_4[16] <= 128'h0F8001F0000000000000000000000000;
                          char22_4[17] <= 128'h1F0001F0000000000000000000000000;
                          char22_4[18] <= 128'h1F0001F0000000000000000000000000;
                          char22_4[19] <= 128'h1F0001F0000000000000000000000000;
                          char22_4[20] <= 128'h1F0001F0000000000000000000000000;
                          char22_4[21] <= 128'h1F0001F0000000000000000000000000;
                          char22_4[22] <= 128'h1F8001F0000000000000000000000000;
                          char22_4[23] <= 128'h1FC001F0000000000000000000000000;
                          char22_4[24] <= 128'h0FC001F0000000000000000000000000;
                          char22_4[25] <= 128'h0FF003E0000000000000000000000000;
                          char22_4[26] <= 128'h07F803C0000000000000000000000000;
                          char22_4[27] <= 128'h03FE0F80000000000000000000000000;
                          char22_4[28] <= 128'h01FF9F00000000000000000000000000;
                          char22_4[29] <= 128'h00FFFE00000000000000000000000000;
                          char22_4[30] <= 128'h003FF800000000000000000000000000;
                          char22_4[31] <= 128'h007FFC00000000000000000000000000;
                          char22_4[32] <= 128'h01F7FF00000000000000000000000000;
                          char22_4[33] <= 128'h03E1FF80000000000000000000000000;
                          char22_4[34] <= 128'h07C07FC0000000000000000000000000;
                          char22_4[35] <= 128'h0F801FE0000000000000000000000000;
                          char22_4[36] <= 128'h0F800FE0000000000000000000000000;
                          char22_4[37] <= 128'h1F0007F0000000000000000000000000;
                          char22_4[38] <= 128'h1F0003F0000000000000000000000000;
                          char22_4[39] <= 128'h3E0001F8000000000000000000000000;
                          char22_4[40] <= 128'h3E0001F8000000000000000000000000;
                          char22_4[41] <= 128'h3E0001F8000000000000000000000000;
                          char22_4[42] <= 128'h3E0000F8000000000000000000000000;
                          char22_4[43] <= 128'h3E0000F8000000000000000000000000;
                          char22_4[44] <= 128'h3E0000F8000000000000000000000000;
                          char22_4[45] <= 128'h3E0000F8000000000000000000000000;
                          char22_4[46] <= 128'h1F0001F0000000000000000000000000;
                          char22_4[47] <= 128'h1F0001F0000000000000000000000000;
                          char22_4[48] <= 128'h0F8003E0000000000000000000000000;
                          char22_4[49] <= 128'h0FC003E0000000000000000000000000;
                          char22_4[50] <= 128'h07E007C0000000000000000000000000;
                          char22_4[51] <= 128'h01F83F80000000000000000000000000;
                          char22_4[52] <= 128'h00FFFE00000000000000000000000000;
                          char22_4[53] <= 128'h003FF800000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//8
                    4'd9: begin
                          char22_4[0] <= 128'h00000000000000000000000000000000;
                          char22_4[1] <= 128'h00000000000000000000000000000000;
                          char22_4[2] <= 128'h00000000000000000000000000000000;
                          char22_4[3] <= 128'h00000000000000000000000000000000;
                          char22_4[4] <= 128'h00000000000000000000000000000000;
                          char22_4[5] <= 128'h00000000000000000000000000000000;
                          char22_4[6] <= 128'h00000000000000000000000000000000;
                          char22_4[7] <= 128'h00000000000000000000000000000000;
                          char22_4[8] <= 128'h00000000000000000000000000000000;
                          char22_4[9] <= 128'h00000000000000000000000000000000;
                          char22_4[10] <= 128'h003FF000000000000000000000000000;
                          char22_4[11] <= 128'h00FFFC00000000000000000000000000;
                          char22_4[12] <= 128'h01F83F00000000000000000000000000;
                          char22_4[13] <= 128'h03E01F80000000000000000000000000;
                          char22_4[14] <= 128'h07C00F80000000000000000000000000;
                          char22_4[15] <= 128'h0FC007C0000000000000000000000000;
                          char22_4[16] <= 128'h0F8003E0000000000000000000000000;
                          char22_4[17] <= 128'h1F8003E0000000000000000000000000;
                          char22_4[18] <= 128'h1F0003F0000000000000000000000000;
                          char22_4[19] <= 128'h1F0003F0000000000000000000000000;
                          char22_4[20] <= 128'h3F0001F0000000000000000000000000;
                          char22_4[21] <= 128'h3F0001F0000000000000000000000000;
                          char22_4[22] <= 128'h3F0001F8000000000000000000000000;
                          char22_4[23] <= 128'h3F0001F8000000000000000000000000;
                          char22_4[24] <= 128'h3F0001F8000000000000000000000000;
                          char22_4[25] <= 128'h3F0001F8000000000000000000000000;
                          char22_4[26] <= 128'h3F0001F8000000000000000000000000;
                          char22_4[27] <= 128'h3F0001F8000000000000000000000000;
                          char22_4[28] <= 128'h3F0003F8000000000000000000000000;
                          char22_4[29] <= 128'h1F8003F8000000000000000000000000;
                          char22_4[30] <= 128'h1F8007F8000000000000000000000000;
                          char22_4[31] <= 128'h1F800FF8000000000000000000000000;
                          char22_4[32] <= 128'h0FC01FF8000000000000000000000000;
                          char22_4[33] <= 128'h0FE03FF8000000000000000000000000;
                          char22_4[34] <= 128'h07F8FDF8000000000000000000000000;
                          char22_4[35] <= 128'h03FFF9F8000000000000000000000000;
                          char22_4[36] <= 128'h01FFF1F8000000000000000000000000;
                          char22_4[37] <= 128'h003F83F8000000000000000000000000;
                          char22_4[38] <= 128'h000003F0000000000000000000000000;
                          char22_4[39] <= 128'h000003F0000000000000000000000000;
                          char22_4[40] <= 128'h000003F0000000000000000000000000;
                          char22_4[41] <= 128'h000003F0000000000000000000000000;
                          char22_4[42] <= 128'h000007E0000000000000000000000000;
                          char22_4[43] <= 128'h000007E0000000000000000000000000;
                          char22_4[44] <= 128'h000007C0000000000000000000000000;
                          char22_4[45] <= 128'h03C007C0000000000000000000000000;
                          char22_4[46] <= 128'h07C00F80000000000000000000000000;
                          char22_4[47] <= 128'h0FE00F80000000000000000000000000;
                          char22_4[48] <= 128'h0FE01F00000000000000000000000000;
                          char22_4[49] <= 128'h0FE03E00000000000000000000000000;
                          char22_4[50] <= 128'h07E07E00000000000000000000000000;
                          char22_4[51] <= 128'h07F1F800000000000000000000000000;
                          char22_4[52] <= 128'h03FFF000000000000000000000000000;
                          char22_4[53] <= 128'h00FFC000000000000000000000000000;
                          char22_4[54] <= 128'h00000000000000000000000000000000;
                          char22_4[55] <= 128'h00000000000000000000000000000000;
                          char22_4[56] <= 128'h00000000000000000000000000000000;
                          char22_4[57] <= 128'h00000000000000000000000000000000;
                          char22_4[58] <= 128'h00000000000000000000000000000000;
                          char22_4[59] <= 128'h00000000000000000000000000000000;
                          char22_4[60] <= 128'h00000000000000000000000000000000;
                          char22_4[61] <= 128'h00000000000000000000000000000000;
                          char22_4[62] <= 128'h00000000000000000000000000000000;
                          char22_4[63] <= 128'h00000000000000000000000000000000;
                    end//9
                    default: begin
                        char22_4[0] <= char22_4[0];
                        char22_4[1] <= char22_4[1];
                        char22_4[2] <= char22_4[2];
                        char22_4[3] <= char22_4[3];
                        char22_4[4] <= char22_4[4];
                        char22_4[5] <= char22_4[5];
                        char22_4[6] <= char22_4[6];
                        char22_4[7] <= char22_4[7];
                        char22_4[8] <= char22_4[8];
                        char22_4[9] <= char22_4[9];
                        char22_4[10] <= char22_4[10];
                        char22_4[11] <= char22_4[11];
                        char22_4[12] <= char22_4[12];
                        char22_4[13] <= char22_4[13];
                        char22_4[14] <= char22_4[14];
                        char22_4[15] <= char22_4[15];
                        char22_4[16] <= char22_4[16];
                        char22_4[17] <= char22_4[17];
                        char22_4[18] <= char22_4[18];
                        char22_4[19] <= char22_4[19];
                        char22_4[20] <= char22_4[20];
                        char22_4[21] <= char22_4[21];
                        char22_4[22] <= char22_4[22];
                        char22_4[23] <= char22_4[23];
                        char22_4[24] <= char22_4[24];
                        char22_4[25] <= char22_4[25];
                        char22_4[26] <= char22_4[26];
                        char22_4[27] <= char22_4[27];
                        char22_4[28] <= char22_4[28];
                        char22_4[29] <= char22_4[29];
                        char22_4[30] <= char22_4[30];
                        char22_4[31] <= char22_4[31];
                        char22_4[32] <= char22_4[32];
                        char22_4[33] <= char22_4[33];
                        char22_4[34] <= char22_4[34];
                        char22_4[35] <= char22_4[35];
                        char22_4[36] <= char22_4[36];
                        char22_4[37] <= char22_4[37];
                        char22_4[38] <= char22_4[38];
                        char22_4[39] <= char22_4[39];
                        char22_4[40] <= char22_4[40];
                        char22_4[41] <= char22_4[41];
                        char22_4[42] <= char22_4[42];
                        char22_4[43] <= char22_4[43];
                        char22_4[44] <= char22_4[44];
                        char22_4[45] <= char22_4[45];
                        char22_4[46] <= char22_4[46];
                        char22_4[47] <= char22_4[47];
                        char22_4[48] <= char22_4[48];
                        char22_4[49] <= char22_4[49];
                        char22_4[50] <= char22_4[50];
                        char22_4[51] <= char22_4[51];
                        char22_4[52] <= char22_4[52];
                        char22_4[53] <= char22_4[53];
                        char22_4[54] <= char22_4[54];
                        char22_4[55] <= char22_4[55];
                        char22_4[56] <= char22_4[56];
                        char22_4[57] <= char22_4[57];
                        char22_4[58] <= char22_4[58];
                        char22_4[59] <= char22_4[59];
                        char22_4[60] <= char22_4[60];
                        char22_4[61] <= char22_4[61];
                        char22_4[62] <= char22_4[62];
                        char22_4[63] <= char22_4[63];
                    end
                endcase
        
    
  
  
 char22_3[0] <= 32'h00000000;
 char22_3[1] <= 32'h00000000;
 char22_3[2] <= 32'h00000000;
 char22_3[3] <= 32'h00000000;
 char22_3[4] <= 32'h00000000;
 char22_3[5] <= 32'h00000000;
 char22_3[6] <= 32'h00000000;
 char22_3[7] <= 32'h00000000;
 char22_3[8] <= 32'h00000000;
 char22_3[9] <= 32'h00000000;
 char22_3[10] <= 32'h00000000;
 char22_3[11] <= 32'h00000000;
 char22_3[12] <= 32'h00000000;
 char22_3[13] <= 32'h00000000;
 char22_3[14] <= 32'h00000000;
 char22_3[15] <= 32'h00000000;
 char22_3[16] <= 32'h00000000;
 char22_3[17] <= 32'h00000000;
 char22_3[18] <= 32'h00000000;
 char22_3[19] <= 32'h00000000;
 char22_3[20] <= 32'h00000000;
 char22_3[21] <= 32'h00000000;
 char22_3[22] <= 32'h00000000;
 char22_3[23] <= 32'h00000000;
 char22_3[24] <= 32'h00000000;
 char22_3[25] <= 32'h00000000;
 char22_3[26] <= 32'h00000000;
 char22_3[27] <= 32'h00000000;
 char22_3[28] <= 32'h00000000;
 char22_3[29] <= 32'h00000000;
 char22_3[30] <= 32'h00000000;
 char22_3[31] <= 32'h00000000;
 char22_3[32] <= 32'h00000000;
 char22_3[33] <= 32'h00000000;
 char22_3[34] <= 32'h00000000;
 char22_3[35] <= 32'h00000000;
 char22_3[36] <= 32'h00000000;
 char22_3[37] <= 32'h00000000;
 char22_3[38] <= 32'h00000000;
 char22_3[39] <= 32'h00000000;
 char22_3[40] <= 32'h00000000;
 char22_3[41] <= 32'h00000000;
 char22_3[42] <= 32'h00000000;
 char22_3[43] <= 32'h00000000;
 char22_3[44] <= 32'h00000000;
 char22_3[45] <= 32'h00000000;
 char22_3[46] <= 32'h07E00000;
 char22_3[47] <= 32'h0FF00000;
 char22_3[48] <= 32'h0FF00000;
 char22_3[49] <= 32'h0FF00000;
 char22_3[50] <= 32'h0FF00000;
 char22_3[51] <= 32'h0FF00000;
 char22_3[52] <= 32'h0FF00000;
 char22_3[53] <= 32'h07E00000;
 char22_3[54] <= 32'h00000000;
 char22_3[55] <= 32'h00000000;
 char22_3[56] <= 32'h00000000;
 char22_3[57] <= 32'h00000000;
 char22_3[58] <= 32'h00000000;
 char22_3[59] <= 32'h00000000;
 char22_3[60] <= 32'h00000000;
 char22_3[61] <= 32'h00000000;
 char22_3[62] <= 32'h00000000;
 char22_3[63] <= 32'h00000000;
 
 

 
 char[  0] <= {char00[0],char0[0]};
 char[  1] <= {char00[1],char0[1]};
 char[  2] <= {char00[2],char0[2]};
 char[  3] <= {char00[3],char0[3]};
 char[  4] <= {char00[4],char0[4]};
 char[  5] <= {char00[5],char0[5]};
 char[  6] <= {char00[6],char0[6]};
 char[  7] <= {char00[7],char0[7]};
 char[  8] <= {char00[8],char0[8]};
 char[  9] <= {char00[9],char0[9]};
 char[10] <= {char00[10],char0[10]};
 char[11] <= {char00[11],char0[11]};
 char[12] <= {char00[12],char0[12]};
 char[13] <= {char00[13],char0[13]};
 char[14] <= {char00[14],char0[14]};
 char[15] <= {char00[15],char0[15]};
 char[16] <= {char00[16],char0[16]};
 char[17] <= {char00[17],char0[17]};
 char[18] <= {char00[18],char0[18]};
 char[19] <= {char00[19],char0[19]};
 char[20] <= {char00[20],char0[20]};
 char[21] <= {char00[21],char0[21]};
 char[22] <= {char00[22],char0[22]};
 char[23] <= {char00[23],char0[23]};
 char[24] <= {char00[24],char0[24]};
 char[25] <= {char00[25],char0[25]};
 char[26] <= {char00[26],char0[26]};
 char[27] <= {char00[27],char0[27]};
 char[28] <= {char00[28],char0[28]};
 char[29] <= {char00[29],char0[29]};
 char[30] <= {char00[30],char0[30]};
 char[31] <= {char00[31],char0[31]};
 char[32] <= {char00[32],char0[32]};
 char[33] <= {char00[33],char0[33]};
 char[34] <= {char00[34],char0[34]};
 char[35] <= {char00[35],char0[35]};
 char[36] <= {char00[36],char0[36]};
 char[37] <= {char00[37],char0[37]};
 char[38] <= {char00[38],char0[38]};
 char[39] <= {char00[39],char0[39]};
 char[40] <= {char00[40],char0[40]};
 char[41] <= {char00[41],char0[41]};
 char[42] <= {char00[42],char0[42]};
 char[43] <= {char00[43],char0[43]};
 char[44] <= {char00[44],char0[44]};
 char[45] <= {char00[45],char0[45]};
 char[46] <= {char00[46],char0[46]};
 char[47] <= {char00[47],char0[47]};
 char[48] <= {char00[48],char0[48]};
 char[49] <= {char00[49],char0[49]};
 char[50] <= {char00[50],char0[50]};
 char[51] <= {char00[51],char0[51]};
 char[52] <= {char00[52],char0[52]};
 char[53] <= {char00[53],char0[53]};
 char[54] <= {char00[54],char0[54]};
 char[55] <= {char00[55],char0[55]};
 char[56] <= {char00[56],char0[56]};
 char[57] <= {char00[57],char0[57]};
 char[58] <= {char00[58],char0[58]};
 char[59] <= {char00[59],char0[59]};
 char[60] <= {char00[60],char0[60]};
 char[61] <= {char00[61],char0[61]};
 char[62] <= {char00[62],char0[62]};
 char[63] <= {char00[63],char0[63]};
 char[64] <= {char11[0],char1[0]};
 char[65] <= {char11[1],char1[1]};
 char[66] <= {char11[2],char1[2]};
 char[67] <= {char11[3],char1[3]};
 char[68] <= {char11[4],char1[4]};
 char[69] <= {char11[5],char1[5]};
 char[70] <= {char11[6],char1[6]};
 char[71] <= {char11[7],char1[7]};
 char[72] <= {char11[8],char1[8]};
 char[73] <= {char11[9],char1[9]};
 char[74] <= {char11[10],char1[10]};
 char[75] <= {char11[11],char1[11]};
 char[76] <= {char11[12],char1[12]};
 char[77] <= {char11[13],char1[13]};
 char[78] <= {char11[14],char1[14]};
 char[79] <= {char11[15],char1[15]};
 char[80] <= {char11[16],char1[16]};
 char[81] <= {char11[17],char1[17]};
 char[82] <= {char11[18],char1[18]};
 char[83] <= {char11[19],char1[19]};
 char[84] <= {char11[20],char1[20]};
 char[85] <= {char11[21],char1[21]};
 char[86] <= {char11[22],char1[22]};
 char[87] <= {char11[23],char1[23]};
 char[88] <= {char11[24],char1[24]};
 char[89] <= {char11[25],char1[25]};
 char[90] <= {char11[26],char1[26]};
 char[91] <= {char11[27],char1[27]};
 char[92] <= {char11[28],char1[28]};
 char[93] <= {char11[29],char1[29]};
 char[94] <= {char11[30],char1[30]};
 char[95] <= {char11[31],char1[31]};
 char[96] <= {char11[32],char1[32]};
 char[97] <= {char11[33],char1[33]};
 char[98] <= {char11[34],char1[34]};
 char[99] <= {char11[35],char1[35]};
 char[100] <= {char11[36],char1[36]};
 char[101] <= {char11[37],char1[37]};
 char[102] <= {char11[38],char1[38]};
 char[103] <= {char11[39],char1[39]};
 char[104] <= {char11[40],char1[40]};
 char[105] <= {char11[41],char1[41]};
 char[106] <= {char11[42],char1[42]};
 char[107] <= {char11[43],char1[43]};
 char[108] <= {char11[44],char1[44]};
 char[109] <= {char11[45],char1[45]};
 char[110] <= {char11[46],char1[46]};
 char[111] <= {char11[47],char1[47]};
 char[112] <= {char11[48],char1[48]};
 char[113] <= {char11[49],char1[49]};
 char[114] <= {char11[50],char1[50]};
 char[115] <= {char11[51],char1[51]};
 char[116] <= {char11[52],char1[52]};
 char[117] <= {char11[53],char1[53]};
 char[118] <= {char11[54],char1[54]};
 char[119] <= {char11[55],char1[55]};
 char[120] <= {char11[56],char1[56]};
 char[121] <= {char11[57],char1[57]};
 char[122] <= {char11[58],char1[58]};
 char[123] <= {char11[59],char1[59]};
 char[124] <= {char11[60],char1[60]};
 char[125] <= {char11[61],char1[61]};
 char[126] <= {char11[62],char1[62]};
 char[127] <= {char11[63],char1[63]};
 
     char[128] <= {char22_0[0],char22_1[0],char22_2[0],char22_3[0],char22_4[0],char2[0]};
     char[129] <= {char22_0[1],char22_1[1],char22_2[1],char22_3[1],char22_4[1],char2[1]};
     char[130] <= {char22_0[2],char22_1[2],char22_2[2],char22_3[2],char22_4[2],char2[2]};
     char[131] <= {char22_0[3],char22_1[3],char22_2[3],char22_3[3],char22_4[3],char2[3]};
     char[132] <= {char22_0[4],char22_1[4],char22_2[4],char22_3[4],char22_4[4],char2[4]};
     char[133] <= {char22_0[5],char22_1[5],char22_2[5],char22_3[5],char22_4[5],char2[5]};
     char[134] <= {char22_0[6],char22_1[6],char22_2[6],char22_3[6],char22_4[6],char2[6]};
     char[135] <= {char22_0[7],char22_1[7],char22_2[7],char22_3[7],char22_4[7],char2[7]};
     char[136] <= {char22_0[8],char22_1[8],char22_2[8],char22_3[8],char22_4[8],char2[8]};
     char[137] <= {char22_0[9],char22_1[9],char22_2[9],char22_3[9],char22_4[9],char2[9]};
     char[138] <= {char22_0[10],char22_1[10],char22_2[10],char22_3[10],char22_4[10],char2[10]};
     char[139] <= {char22_0[11],char22_1[11],char22_2[11],char22_3[11],char22_4[11],char2[11]};
     char[140] <= {char22_0[12],char22_1[12],char22_2[12],char22_3[12],char22_4[12],char2[12]};
     char[141] <= {char22_0[13],char22_1[13],char22_2[13],char22_3[13],char22_4[13],char2[13]};
     char[142] <= {char22_0[14],char22_1[14],char22_2[14],char22_3[14],char22_4[14],char2[14]};
     char[143] <= {char22_0[15],char22_1[15],char22_2[15],char22_3[15],char22_4[15],char2[15]};
     char[144] <= {char22_0[16],char22_1[16],char22_2[16],char22_3[16],char22_4[16],char2[16]};
     char[145] <= {char22_0[17],char22_1[17],char22_2[17],char22_3[17],char22_4[17],char2[17]};
     char[146] <= {char22_0[18],char22_1[18],char22_2[18],char22_3[18],char22_4[18],char2[18]};
     char[147] <= {char22_0[19],char22_1[19],char22_2[19],char22_3[19],char22_4[19],char2[19]};
     char[148] <= {char22_0[20],char22_1[20],char22_2[20],char22_3[20],char22_4[20],char2[20]};
     char[149] <= {char22_0[21],char22_1[21],char22_2[21],char22_3[21],char22_4[21],char2[21]};
     char[150] <= {char22_0[22],char22_1[22],char22_2[22],char22_3[22],char22_4[22],char2[22]};
     char[151] <= {char22_0[23],char22_1[23],char22_2[23],char22_3[23],char22_4[23],char2[23]};
     char[152] <= {char22_0[24],char22_1[24],char22_2[24],char22_3[24],char22_4[24],char2[24]};
     char[153] <= {char22_0[25],char22_1[25],char22_2[25],char22_3[25],char22_4[25],char2[25]};
     char[154] <= {char22_0[26],char22_1[26],char22_2[26],char22_3[26],char22_4[26],char2[26]};
     char[155] <= {char22_0[27],char22_1[27],char22_2[27],char22_3[27],char22_4[27],char2[27]};
     char[156] <= {char22_0[28],char22_1[28],char22_2[28],char22_3[28],char22_4[28],char2[28]};
     char[157] <= {char22_0[29],char22_1[29],char22_2[29],char22_3[29],char22_4[29],char2[29]};
     char[158] <= {char22_0[30],char22_1[30],char22_2[30],char22_3[30],char22_4[30],char2[30]};
     char[159] <= {char22_0[31],char22_1[31],char22_2[31],char22_3[31],char22_4[31],char2[31]};
     char[160] <= {char22_0[32],char22_1[32],char22_2[32],char22_3[32],char22_4[32],char2[32]};
     char[161] <= {char22_0[33],char22_1[33],char22_2[33],char22_3[33],char22_4[33],char2[33]};
     char[162] <= {char22_0[34],char22_1[34],char22_2[34],char22_3[34],char22_4[34],char2[34]};
     char[163] <= {char22_0[35],char22_1[35],char22_2[35],char22_3[35],char22_4[35],char2[35]};
     char[164] <= {char22_0[36],char22_1[36],char22_2[36],char22_3[36],char22_4[36],char2[36]};
     char[165] <= {char22_0[37],char22_1[37],char22_2[37],char22_3[37],char22_4[37],char2[37]};
     char[166] <= {char22_0[38],char22_1[38],char22_2[38],char22_3[38],char22_4[38],char2[38]};
     char[167] <= {char22_0[39],char22_1[39],char22_2[39],char22_3[39],char22_4[39],char2[39]};
     char[168] <= {char22_0[40],char22_1[40],char22_2[40],char22_3[40],char22_4[40],char2[40]};
     char[169] <= {char22_0[41],char22_1[41],char22_2[41],char22_3[41],char22_4[41],char2[41]};
     char[170] <= {char22_0[42],char22_1[42],char22_2[42],char22_3[42],char22_4[42],char2[42]};
     char[171] <= {char22_0[43],char22_1[43],char22_2[43],char22_3[43],char22_4[43],char2[43]};
     char[172] <= {char22_0[44],char22_1[44],char22_2[44],char22_3[44],char22_4[44],char2[44]};
     char[173] <= {char22_0[45],char22_1[45],char22_2[45],char22_3[45],char22_4[45],char2[45]};
     char[174] <= {char22_0[46],char22_1[46],char22_2[46],char22_3[46],char22_4[46],char2[46]};
     char[175] <= {char22_0[47],char22_1[47],char22_2[47],char22_3[47],char22_4[47],char2[47]};
     char[176] <= {char22_0[48],char22_1[48],char22_2[48],char22_3[48],char22_4[48],char2[48]};
     char[177] <= {char22_0[49],char22_1[49],char22_2[49],char22_3[49],char22_4[49],char2[49]};
     char[178] <= {char22_0[50],char22_1[50],char22_2[50],char22_3[50],char22_4[50],char2[50]};
     char[179] <= {char22_0[51],char22_1[51],char22_2[51],char22_3[51],char22_4[51],char2[51]};
     char[180] <= {char22_0[52],char22_1[52],char22_2[52],char22_3[52],char22_4[52],char2[52]};
     char[181] <= {char22_0[53],char22_1[53],char22_2[53],char22_3[53],char22_4[53],char2[53]};
     char[182] <= {char22_0[54],char22_1[54],char22_2[54],char22_3[54],char22_4[54],char2[54]};
     char[183] <= {char22_0[55],char22_1[55],char22_2[55],char22_3[55],char22_4[55],char2[55]};
     char[184] <= {char22_0[56],char22_1[56],char22_2[56],char22_3[56],char22_4[56],char2[56]};
     char[185] <= {char22_0[57],char22_1[57],char22_2[57],char22_3[57],char22_4[57],char2[57]};
     char[186] <= {char22_0[58],char22_1[58],char22_2[58],char22_3[58],char22_4[58],char2[58]};
     char[187] <= {char22_0[59],char22_1[59],char22_2[59],char22_3[59],char22_4[59],char2[59]};
     char[188] <= {char22_0[60],char22_1[60],char22_2[60],char22_3[60],char22_4[60],char2[60]};
     char[189] <= {char22_0[61],char22_1[61],char22_2[61],char22_3[61],char22_4[61],char2[61]};
     char[190] <= {char22_0[62],char22_1[62],char22_2[62],char22_3[62],char22_4[62],char2[62]};
     char[191] <= {char22_0[63],char22_1[63],char22_2[63],char22_3[63],char22_4[63],char2[63]};

 char[192] <= 512'h0;
     char[193] <= 512'h0;
     char[194] <= 512'h0;
     char[195] <= 512'h0;
     char[196] <= 512'h0;
     char[197] <= 512'h0;
     char[198] <= 512'h0;
     char[199] <= 512'h0;
     char[200] <= 512'h0;
     char[201] <= 512'h0;
     char[202] <= 512'h0;
     char[203] <= 512'h0;
     char[204] <= 512'h0;
     char[205] <= 512'h0;
     char[206] <= 512'h0;
     char[207] <= 512'h0;
     char[208] <= 512'h0;
     char[209] <= 512'h0;
     char[210] <= 512'h0;
     char[211] <= 512'h0;
     char[212] <= 512'h0;
     char[213] <= 512'h0;
     char[214] <= 512'h0;
     char[215] <= 512'h0;
     char[216] <= 512'h0;
     char[217] <= 512'h0;
     char[218] <= 512'h0;
     char[219] <= 512'h0;
     char[220] <= 512'h0;
     char[221] <= 512'h0;
     char[222] <= 512'h0;
     char[223] <= 512'h0;
     char[224] <= 512'h0;
     char[225] <= 512'h0;
     char[226] <= 512'h0;
     char[227] <= 512'h0;
     char[228] <= 512'h0;
     char[229] <= 512'h0;
     char[230] <= 512'h0;
     char[231] <= 512'h0;
     char[232] <= 512'h0;
     char[233] <= 512'h0;
     char[234] <= 512'h0;
     char[235] <= 512'h0;
     char[236] <= 512'h0;
     char[237] <= 512'h0;
     char[238] <= 512'h0;
     char[239] <= 512'h0;
     char[240] <= 512'h0;
     char[241] <= 512'h0;
     char[242] <= 512'h0;
     char[243] <= 512'h0;
     char[244] <= 512'h0;
     char[245] <= 512'h0;
     char[246] <= 512'h0;
     char[247] <= 512'h0;
     char[248] <= 512'h0;
     char[249] <= 512'h0;
     char[250] <= 512'h0;
     char[251] <= 512'h0;
     char[252] <= 512'h0;
     char[253] <= 512'h0;
     char[254] <= 512'h0;
     char[255] <= 512'h0;
     char[256] <= 512'h0;
     char[257] <= 512'h0;
     char[258] <= 512'h0;
     char[259] <= 512'h0;
     char[260] <= 512'h0;
     char[261] <= 512'h0;
     char[262] <= 512'h0;
     char[263] <= 512'h0;
     char[264] <= 512'h0;
     char[265] <= 512'h0;
     char[266] <= 512'h0;
     char[267] <= 512'h0;
     char[268] <= 512'h0;
     char[269] <= 512'h0;
     char[270] <= 512'h0;
     char[271] <= 512'h0;
     char[272] <= 512'h0;
     char[273] <= 512'h0;
     char[274] <= 512'h0;
     char[275] <= 512'h0;
     char[276] <= 512'h0;
     char[277] <= 512'h0;
     char[278] <= 512'h0;
     char[279] <= 512'h0;
     char[280] <= 512'h0;
     char[281] <= 512'h0;
     char[282] <= 512'h0;
     char[283] <= 512'h0;
     char[284] <= 512'h0;
     char[285] <= 512'h0;
     char[286] <= 512'h0;
     char[287] <= 512'h0;
     char[288] <= 512'h0;
     char[289] <= 512'h0;
     char[290] <= 512'h0;
     char[291] <= 512'h0;
     char[292] <= 512'h0;
     char[293] <= 512'h0;
     char[294] <= 512'h0;
     char[295] <= 512'h0;
     char[296] <= 512'h0;
     char[297] <= 512'h0;
     char[298] <= 512'h0;
     char[299] <= 512'h0;
     char[300] <= 512'h0;
     char[301] <= 512'h0;
     char[302] <= 512'h0;
     char[303] <= 512'h0;
     char[304] <= 512'h0;
     char[305] <= 512'h0;
     char[306] <= 512'h0;
     char[307] <= 512'h0;
     char[308] <= 512'h0;
     char[309] <= 512'h0;
     char[310] <= 512'h0;
     char[311] <= 512'h0;
     char[312] <= 512'h0;
     char[313] <= 512'h0;
     char[314] <= 512'h0;
     char[315] <= 512'h0;
     char[316] <= 512'h0;
     char[317] <= 512'h0;
     char[318] <= 512'h0;
     char[319] <= 512'h0;
     char[320] <= 512'h0;
     char[321] <= 512'h0;
     char[322] <= 512'h0;
     char[323] <= 512'h0;
     char[324] <= 512'h0;
     char[325] <= 512'h0;
     char[326] <= 512'h0;
     char[327] <= 512'h0;
     char[328] <= 512'h0;
     char[329] <= 512'h0;
     char[330] <= 512'h0;
     char[331] <= 512'h0;
     char[332] <= 512'h0;
     char[333] <= 512'h0;
     char[334] <= 512'h0;
     char[335] <= 512'h0;
     char[336] <= 512'h0;
     char[337] <= 512'h0;
     char[338] <= 512'h0;
     char[339] <= 512'h0;
     char[340] <= 512'h0;
     char[341] <= 512'h0;
     char[342] <= 512'h0;
     char[343] <= 512'h0;
     char[344] <= 512'h0;
     char[345] <= 512'h0;
     char[346] <= 512'h0;
     char[347] <= 512'h0;
     char[348] <= 512'h0;
     char[349] <= 512'h0;
     char[350] <= 512'h0;
     char[351] <= 512'h0;
     char[352] <= 512'h0;
     char[353] <= 512'h0;
     char[354] <= 512'h0;
     char[355] <= 512'h0;
     char[356] <= 512'h0;
     char[357] <= 512'h0;
     char[358] <= 512'h0;
     char[359] <= 512'h0;
     char[360] <= 512'h0;
     char[361] <= 512'h0;
     char[362] <= 512'h0;
     char[363] <= 512'h0;
     char[364] <= 512'h0;
     char[365] <= 512'h0;
     char[366] <= 512'h0;
     char[367] <= 512'h0;
     char[368] <= 512'h0;
     char[369] <= 512'h0;
     char[370] <= 512'h0;
     char[371] <= 512'h0;
     char[372] <= 512'h0;
     char[373] <= 512'h0;
     char[374] <= 512'h0;
     char[375] <= 512'h0;
     char[376] <= 512'h0;
     char[377] <= 512'h0;
     char[378] <= 512'h0;
     char[379] <= 512'h0;
     char[380] <= 512'h0;
     char[381] <= 512'h0;
     char[382] <= 512'h0;
     char[383] <= 512'h0;
     char[384] <= 512'h0;
     char[385] <= 512'h0;
     char[386] <= 512'h0;
     char[387] <= 512'h0;
     char[388] <= 512'h0;
     char[389] <= 512'h0;
     char[390] <= 512'h0;
     char[391] <= 512'h0;
     char[392] <= 512'h0;
     char[393] <= 512'h0;
     char[394] <= 512'h0;
     char[395] <= 512'h0;
     char[396] <= 512'h0;
     char[397] <= 512'h0;
     char[398] <= 512'h0;
     char[399] <= 512'h0;
     char[400] <= 512'h0;
     char[401] <= 512'h0;
     char[402] <= 512'h0;
     char[403] <= 512'h0;
     char[404] <= 512'h0;
     char[405] <= 512'h0;
     char[406] <= 512'h0;
     char[407] <= 512'h0;
     char[408] <= 512'h0;
     char[409] <= 512'h0;
     char[410] <= 512'h0;
     char[411] <= 512'h0;
     char[412] <= 512'h0;
     char[413] <= 512'h0;
     char[414] <= 512'h0;
     char[415] <= 512'h0;
     char[416] <= 512'h0;
     char[417] <= 512'h0;
     char[418] <= 512'h0;
     char[419] <= 512'h0;
     char[420] <= 512'h0;
     char[421] <= 512'h0;
     char[422] <= 512'h0;
     char[423] <= 512'h0;
     char[424] <= 512'h0;
     char[425] <= 512'h0;
     char[426] <= 512'h0;
     char[427] <= 512'h0;
     char[428] <= 512'h0;
     char[429] <= 512'h0;
     char[430] <= 512'h0;
     char[431] <= 512'h0;
     char[432] <= 512'h0;
     char[433] <= 512'h0;
     char[434] <= 512'h0;
     char[435] <= 512'h0;
     char[436] <= 512'h0;
     char[437] <= 512'h0;
     char[438] <= 512'h0;
     char[439] <= 512'h0;
     char[440] <= 512'h0;
     char[441] <= 512'h0;
     char[442] <= 512'h0;
     char[443] <= 512'h0;
     char[444] <= 512'h0;
     char[445] <= 512'h0;
     char[446] <= 512'h0;
     char[447] <= 512'h0;
     char[448] <= 512'h0;
     char[449] <= 512'h0;
     char[450] <= 512'h0;
     char[451] <= 512'h0;
     char[452] <= 512'h0;
     char[453] <= 512'h0;
     char[454] <= 512'h0;
     char[455] <= 512'h0;
     char[456] <= 512'h0;
     char[457] <= 512'h0;
     char[458] <= 512'h0;
     char[459] <= 512'h0;
     char[460] <= 512'h0;
     char[461] <= 512'h0;
     char[462] <= 512'h0;
     char[463] <= 512'h0;
     char[464] <= 512'h0;
     char[465] <= 512'h0;
     char[466] <= 512'h0;
     char[467] <= 512'h0;
     char[468] <= 512'h0;
     char[469] <= 512'h0;
     char[470] <= 512'h0;
     char[471] <= 512'h0;
     char[472] <= 512'h0;
     char[473] <= 512'h0;
     char[474] <= 512'h0;
     char[475] <= 512'h0;
     char[476] <= 512'h0;
     char[477] <= 512'h0;
     char[478] <= 512'h0;
     char[479] <= 512'h0;
end

always @(posedge vga_clk , posedge sys_rst) begin
     if(sys_rst)begin
        pix_data <=black;
     end
     else if (pix_x<512 && char[pix_y][10'd255-pix_x] == 1'b1)
        /*if (pix_x >=416 && pix_y >= 128) pix_data <= white;
        else */pix_data <=blue;
     else
        pix_data <=white;
     
        
end

endmodule

module vga(//clk ��25MHZ
input wire sys_clk,
input wire sys_rst,
input wire[3:0] stat,
input wire [2:0]swi,

output wire hsync,
output wire vsync,
output wire [11:0]vga_rgb
);
wire [9:0] pix_x;
wire [9:0] pix_y;
wire [11:0] pix_data;
wire clk_25m;
vga_control vc(
clk_25m ,  sys_rst ,  pix_data  ,  pix_x  , pix_y  , hsync,  vsync  ,  vga_rgb   
);
vga_draw vd(clk_25m , sys_rst , stat , swi  ,  pix_x , pix_y , pix_data );
Get25Clk Gc(sys_clk  ,sys_rst ,clk_25m);
endmodule

module Get25Clk(input sys_clk,input rst,output reg clk_25m);//��Ƶ��

parameter period =4;
reg[3:0] cnt;
always@(posedge sys_clk,posedge rst )begin
    if(rst)begin
        cnt<=0;
        clk_25m<=0;
        end
     else
           if(cnt==((period>>1)-1)) begin
           clk_25m <=~clk_25m;
           cnt<= 0;
           end 
           else begin
            cnt<=cnt+1;
            end
     end
endmodule
